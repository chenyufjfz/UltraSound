��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��։�������7��*`�ԇ��h��U
�~�a�������.H��N��Y9Ύ�2��3�MT�������-8]#�X̵���lV``�^��k(C6˞��w��7�w�T]U:⡇J?��\f�խ�@��R@���>I6�Y���٦��bQ�ayڼH�������u"�G�Jn/0k�؆-1k;�!��� ƀg Y�ƳA¹�1&t����C@�!Q�p,婕��'��^F"`�'�ar��FRօ6��!Kx!@c�V`�HjR��BBG�_	 �,8�6R>(?�=]=���{۝s�H���'�c !ΐ/��A*�/��~D KmgH�~:�?I���9� ;b1�D���an��˅�E����_G'�`-��s����Ũ���)�dtE��� e�ä
zS�Br��` )��j�흿c
z�7��1� ]�����8kQT3�Q�Qm+��%]�
Sp�	[6�*�9�ϐ��c�0��8�<!�T�(�~�Â�57y�5�"0�Pl�eg9�Ӯ[�1���]`D���쒦]�l���i � ����)F{�`��G�k��j�r�
���C��%e/�ڝ�J2�f=�D�%�h�q@�iG�������p)�����
lO��bc��P�o��xr��&��HI�����:�`���W�F���fk���d>�k�a��I�Ο#�(&u��EM����6���y���r��؄��G�}^0�k���o�^Z��&v	MMJ֮�] M5���n����xJ�ȃ����c%%��y�QYH�ܵm����Ҫ�>��/�
tZRT��-ya�C^�_s�Y�u�!WSW���:�}V����k��¹3gU��GX{e��|n)vp��6�Q�`>��Ո-B�xӵ��w�+�S �7��&*�y�~�(�%���A��VL:j�_�h7�b�ꚾPF]�D�ȷ���8!�%R�:���*��M,����&?�F��P�?Z�4EVȎ�:�0ڢ�%J�Dz)P�C�$��;yK ,�������0ʰ�i�ƺ�%�:���V�^�2Է��3<}����՘����~g؟��� g��y����BHֺ�.�]�/5Ydi��oI���@ݓ����х@=:��l�0��Ó��t%�cDJ#�9^��̎����c<�I,�L� �'B���G=�;��ҙ�)�K�$$dR&��h�y�4�Қ�Kh�j�4@���M���!�û@�2:��ۓ��2���u4�-�f�e�1@�-hB��)��]��kX:��ڮİ���Ʈ�j{eK.qx�ix�Y�jz܌O��,��b�����-��"�aR�Fh� 7�Ly�<�R_�ia���]HH|��-5!=�|i��-���y���b|�r��\��ě*M��e�1�0�jr�!Ki�d@��Gd#��T\K�U���,�@?���k�^�o��+VÆ��k⚾�{!�X��!g�ȣ��pb�6g��}|�غ�����6�Ƶ�MI���X�X��[���u��o�Bk����a�a�֎N���ʿ������1�OG�	�q�v,�[�����ؠ��RZIb��NP�?����Ƥ�r�xx��G�/b�J%{�$g"?��NVw��F=�DDj��:/�3e�I�x��PP�0Q���g����2����lׇ�]�E�4`�>����d���m(�Wdϋj���5�TK�[cM� �?�çlAAm0,���*�2���E��t=�Jx���e��G��bzs�I4�--�rp��������<XM�Du�p�
D�(7үԍ��+W�_QN"L�X��]p^uU9�6�����jn��H�v^)��e݇8�Gdw�>$]�d���#U�h��$�N�H.�������D8Q�U����� �ȅ	�b�T�x�7W���W�ޝ�^OH�%ѽ����W'��
���F#��/C�j�'tICT�~�Lƚ)��hCj 8�'�&�(Q|�����c��A3D�a�͘�c�6+@����=X�Vb�B2�|�2H*�������H����j���qݬ[�<�Woɭ�L��c�k�Q����Оe�^a��o|^+�uΥ�8�B>��J�]z�X@sx�i����9$~��O�+��2�tn����=�
��@�f���<?�|�y�ܯ�!q;����m+��� �={���'M�3��w��	��ɿ��6f��[�lȕD#s}�}��As奎ĎH'���`��l�)�*$h�-w�f��`�Zq���Q�㨰��6#�+�<x������<cW���c��L�
 Ev:���S�zv+���d�A�P��"C��d\�$­A�1yV3��٠�"9@:����0&Eg�aT�f\�$%%�mPg=^~�h����Nd��<&��BR��i �����a��VE����"� �IWgA��ExtL#Z���A��o{Za@�A�_��h�5J6�:�?���żL�2�D������G��x<I��Ŏ�w�(�	O�+�ϟ�1R<F<,/fC{�Qx��1`bdHBgX�S�����Y�z����t��:��
?+�
��`�]M��3|��Qn|���<�g����s�HI�l���?�uj<Geo�ߡ �##$�F����~�S#4��O�X��to�����f����?�L�O�7����!n�9��)�w^ؾ�\y�[���)LO�� (��=⺲�gٮ�vƑ�.��W�k�����x��Kt�cBx� p�S�@!����q9[�?���[��hG?(���=~�o��)�e%zG���dft{p-��鏺"&��qds�L�w;s�ݟ�k����}#�X�ъ6Wە�1�w�נ�K�B���&j��Q�VE�ը9��R�mRU�sz�@ȵ��Ɔ����gm��n����ٕb-���@���-�׀�{�6��wP"�����Ϩ�6v-{Ar�3��B0)~�}�ց����k�$��,"�'��-L"։�+\�)`E�bؿ� �51��4���j	��bH�v����A[���$�@��`,�a�����xB@��n��ƶ�|��v�z<=2��)8Vœy�z>)��_�Q����!^~h��S�]5�H��,�š�SF���P��&٪���ր�.� �<���k�f�T�`��Յ�d�7�vm\�K�!ok+7��,�T���z���4��읁�G��i%H��-����y��m�=i釨u�iT&�����"`7�fn�_Ef�c��:V���S�L{-�<�o4��˝%K�׃��˜V)�H��u�g�g�d�RHk�Y�,xN������9��O��=�,�|͓�F����DZ�7�֪��1B��Egj�e�:�{p%%�-��Op�A@��K� F1��?��%͝�M��u�om�%%+�ח9r��I/���!�|���xvK��gN�<�)����Q�K%��ً�ND��ͽ+�=}�u��~߱T@Vn��a�����z��n�pWqUӍ��Z���zן�#�㐯��r=5O���.NV�����Ԣ�C�H�V
��9��^���b����%�EEi|��~iP��_�f��R>%��NjXs���El�-�It�a�`<mi
?#���9'�;jN:�M?7@�ݐZ�JN����:�g��XJ�����=���?E�R��ո���ח�����x�G�,���B<���͘Gh$.T[#]K�9�{9z�V�ҸL3U��D�$���953&���|��;��Qٶ�Ӧ�y�AT�0gM��N;nsC*�p37���#mۤ�3��cG�ӥ��Y��jcc��U%8gqq' ā���fk��%T�j(^L>�?aR��3��Z�ge�Kv �l��go��^N̠k�s��	�'4��Ӧ�;(���1���/� �xg�n�}�R����.�q��#�`z9�E]/��u92[oz�y�oJU�o����{� _)��oi�|�鼶T�"�)�6��]�@]gS`�������c�� !�&�Tzk��WZe�WKY�1��B��;� �Tru��T�\V�qC�@�ج>*�U��݈�D��P��d�2�� jAK%�ǒ[H��?vaA�����YN��<����]5��k�����:��_h!�+�����ᚸ�����B����WVW!v?���Ln�����bɥ�0���i)��i��	_���
���ϖk_O�tp�"��>T�Wsy�:(^���
�Ϳ9F(�w�OP��x>��t��f�7?ry�I^Иu-;,l?e̢>;�E�1�xQo��#7���^2&��8m���7:M�-h/�sWl��:m��&����j��'�߈��r��G�8�󫊽@Y��6[����{�: I���̅����QҪ�]x��s(W��j��c�}O�7��۪D
-8�V�hu�p�,�V馜]��w���C��k2��'3H��6�z��M��#̰C�[�g4���O~V6*�;���m5 Z���/"�kq�����&$��t
�r�I+e˕ՔG�0���Ĳ���U�T�3!.&�.�b�G�sxV3�^>���������������f��ݳ�*FD?��n��i��y�\��KO���5��sG�� ��ʚKF2��w�2.q�R_�td���&�`�߶����b9��{�m���UGH��Z٘�S�6@�=�G$%Yz���A]|�QO6߹V)�~��h6yp��qU��v�ٮ�1����ǻ�u��;G��
�a_�پ@�ʣ���닚�ZzWT��I=;�����'R�5H�>���M��+j���i;M�ְG���n5/�9^����Q�?�hiԃÛc����{�z_ƽ,s����\�d�x��X^�L:�j�T8^�%$���w��=��"UN���Ր�!�+R�PN/g���.Cl��m��!R�$S��6X��2��oj4�e�gE�&}�Ѱ���z���s�ė�.�|äHl9��EOk�6��l�l\�n�a]px��P�Y�`���ܼl�?�؋�'�����J�r�
��4�4.��W���n�ݒ��X��2?�P&�=��i`�C��������n�^��_���j��;b ��r��^~"h{,��(��;������B�%�e��H��6�(\��$��`�ⱓi+���'�zFD����ۭ� �~�����m���ɸ)a�>��j�%%zhJ�B���~�T#"0�]+f�(T7�����,�D�E��_ۨo��(�t~םS���Öߊ_��������m�h�*5��l���g1C��b�.�K/��Z�T��N{�٪�c���E�j�,ճ�\��L'],[L3*V7�P�rJ�H�Ch�(PS�r���=���o5���{�p�/���؛����+H��N�jT����N�g�Uk���6 ����R?�����10H
�ur�ݽ�}O}�Ǐ. �U(�#z�]�&ʳ���}8;~�C��X���H�~�]͹\����2�j}�"�>���F�+8����Kᒮ�qq/ד��"��ܽ�}�_�e+���jK�=�M���Ž��`;�-"�9عB?fߊ�6V��/ޮ�}�#j���v3$�ꅥ����H�x��K���H����$R�F�V�j�]p�g\<��1�_��`->�x`�u!��īm��B���*?����M�\�Yޅ4�A�6."G�\ap������;��6��,��6������R���Y�'�S�(u�1��Y���W�P�H"��at�Q�ڙ�D7n�k|B�L�"�K_�DzxJ҉D�Q:�6gyԀ�<�نC>��I(�������dY����Kf�t�;/!Яa?�g��s�է��˞z�2��
&+A��R,� ���9���������P�A��Z][��`̷�[K���b�&�ݒ��{���ƾ�O%l���_��N��:�[GC��U��("�AS�jϟ�R��A����f^ަ��#�^ed�ԥ�@*��k��~�#Z��p������Xq�P{ɕ+�6�3�T����uC;4�wG@gcN��9K�C�� ��,S�� �I#��J��0ઁ�zB�]`�ħ@������nQi�\��LY���[�,�A�����̫���U���f����JY����H�ɺ~��9u��2�q�ZP/�t�Y�E�>�qf�WN2��#Scg� ���w���� �W�R�mA�H�{�� 1��%8�zJP���Ѿyl��ճ�}�$��k�8��MӇ՞��~��R���2�<�6�4�T9c�m��n��Ge>)� ����N5lӵ�~V9~� �� ��u���,%v�ӮPې��&���*����w�o�J�UsA�c{y��>�L ļ{i�W���|�զ!�?@@S�OH$����G+��_�7�.�+��f�-�KǦ����(�aܝ�T�j�T�B�	�&-�\�Tc:֊��*Ì\J3����rs�!ѕ��Z5�X�)��*c��<�J,�(.a{�/ʆ��4�#N�Ep\���m6�W��3��K<S#�^�`�y��28P&(�O�!���z?3�	��+O�>��A��	�T��r6~��$	�B��{�-�T|����n��?]�P--�)��9э�GO�&|�� ��2�,x)_�C7��%����<Ϲz-U~�����|�\����ޏ�V�?���Nkj�K2N<J�p=c_���}��Oj��o~���5.1������d+JQ?��ݪ�4�"F���W�g��id���Y��dt�k`������9�R��ݝ=������f/?؅ˍ�2�`��VGn�y�Wߣ��`��G�Ȧ��4Xz�/X[:h��5�T�"���f`R��vL]@�I���\tZ8B*��Lz�3|���h�>�o�Ӎ�4��hJgT�8�%X�k;.;!^7,;n�G�L��Zn����鉔{�NqƇ
��-/���:t2��qٿ�(;|YO#����c���k6h�J"�w��H��~���r�����B��O:�G��KT�o�!�����o�֘�$�����y���o��B����*2
�}��T���*�`M t�sb���t��D$-N�E�H�A�]�(E7Q]���?�fuGJ�����3{�_�N��f�ٝ{ǩO�{���f�܄z����S36��Ը1o[�
�?���}���X�V)�������CZ������v��n!Ef��᤹L^�������D�bs���YUŉ�0N��"���͐V�˛W[7z�wN��`�������F�\#�	�<<
� oeH�{9���