library verilog;
use verilog.vl_types.all;
entity udp_mac_complete is
    generic(
        REAL_PHY        : integer := 0
    );
    port(
        clk             : in     vl_logic;
        clk_2           : in     vl_logic;
        rst             : in     vl_logic;
        reg_addr        : in     vl_logic_vector(7 downto 0);
        reg_rd          : in     vl_logic;
        reg_wr          : in     vl_logic;
        reg_busy        : out    vl_logic;
        reg_writedata   : in     vl_logic_vector(31 downto 0);
        reg_readdata    : out    vl_logic_vector(31 downto 0);
        tx_clk          : in     vl_logic;
        rx_clk          : in     vl_logic;
        tx_control      : out    vl_logic;
        rx_control      : in     vl_logic;
        rgmii_in        : in     vl_logic_vector(3 downto 0);
        rgmii_out       : out    vl_logic_vector(3 downto 0);
        in_ip_hdr_valid : in     vl_logic;
        in_ip_hdr_ready : out    vl_logic;
        in_ip_dscp      : in     vl_logic_vector(5 downto 0);
        in_ip_ecn       : in     vl_logic_vector(1 downto 0);
        in_ip_length    : in     vl_logic_vector(15 downto 0);
        in_ip_ttl       : in     vl_logic_vector(7 downto 0);
        in_ip_protocol  : in     vl_logic_vector(7 downto 0);
        in_ip_source_ip : in     vl_logic_vector(31 downto 0);
        in_ip_dest_ip   : in     vl_logic_vector(31 downto 0);
        in_ip_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        in_ip_payload_axis_tvalid: in     vl_logic;
        in_ip_payload_axis_tready: out    vl_logic;
        in_ip_payload_axis_tlast: in     vl_logic;
        in_ip_payload_axis_tuser: in     vl_logic;
        tx_udp_hdr_valid: in     vl_logic;
        tx_udp_hdr_ready: out    vl_logic;
        tx_udp_ip_dscp  : in     vl_logic_vector(5 downto 0);
        tx_udp_ip_ecn   : in     vl_logic_vector(1 downto 0);
        tx_udp_ip_ttl   : in     vl_logic_vector(7 downto 0);
        tx_udp_ip_dest_ip: in     vl_logic_vector(31 downto 0);
        tx_udp_source_port: in     vl_logic_vector(15 downto 0);
        tx_udp_dest_port: in     vl_logic_vector(15 downto 0);
        tx_udp_length   : in     vl_logic_vector(15 downto 0);
        tx_udp_checksum : in     vl_logic_vector(15 downto 0);
        tx_udp_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        tx_udp_payload_axis_tvalid: in     vl_logic;
        tx_udp_payload_axis_tready: out    vl_logic;
        tx_udp_payload_axis_tlast: in     vl_logic;
        tx_udp_payload_axis_tuser: in     vl_logic;
        rx_udp_hdr_valid: out    vl_logic;
        rx_udp_hdr_ready: in     vl_logic;
        rx_udp_eth_dest_mac: out    vl_logic_vector(47 downto 0);
        rx_udp_eth_src_mac: out    vl_logic_vector(47 downto 0);
        rx_udp_eth_type : out    vl_logic_vector(15 downto 0);
        rx_udp_ip_version: out    vl_logic_vector(3 downto 0);
        rx_udp_ip_ihl   : out    vl_logic_vector(3 downto 0);
        rx_udp_ip_dscp  : out    vl_logic_vector(5 downto 0);
        rx_udp_ip_ecn   : out    vl_logic_vector(1 downto 0);
        rx_udp_ip_length: out    vl_logic_vector(15 downto 0);
        rx_udp_ip_identification: out    vl_logic_vector(15 downto 0);
        rx_udp_ip_flags : out    vl_logic_vector(2 downto 0);
        rx_udp_ip_fragment_offset: out    vl_logic_vector(12 downto 0);
        rx_udp_ip_ttl   : out    vl_logic_vector(7 downto 0);
        rx_udp_ip_protocol: out    vl_logic_vector(7 downto 0);
        rx_udp_ip_header_checksum: out    vl_logic_vector(15 downto 0);
        rx_udp_ip_source_ip: out    vl_logic_vector(31 downto 0);
        rx_udp_ip_dest_ip: out    vl_logic_vector(31 downto 0);
        rx_udp_source_port: out    vl_logic_vector(15 downto 0);
        rx_udp_dest_port: out    vl_logic_vector(15 downto 0);
        rx_udp_length   : out    vl_logic_vector(15 downto 0);
        rx_udp_checksum : out    vl_logic_vector(15 downto 0);
        rx_udp_payload_axis_tdata: out    vl_logic_vector(7 downto 0);
        rx_udp_payload_axis_tvalid: out    vl_logic;
        rx_udp_payload_axis_tready: in     vl_logic;
        rx_udp_payload_axis_tlast: out    vl_logic;
        rx_udp_payload_axis_tuser: out    vl_logic;
        rx_udp_err      : out    vl_logic;
        local_ip        : out    vl_logic_vector(31 downto 0);
        eth_mode        : out    vl_logic;
        mdc             : out    vl_logic;
        mdio_in         : in     vl_logic;
        mdio_oen        : out    vl_logic;
        mdio_out        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of REAL_PHY : constant is 1;
end udp_mac_complete;
