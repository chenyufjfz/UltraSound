��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�P��9z�7a�U,?�y�"{�Rm�6�¼�L��H�Wl:�j��.����u@X�����b]7u��~V������[Kv�@ъ4gB�䩯ڴO����LHvUmw��[ї:�⻛`CC��;�����@L46�M�p!��ߔ��aP�фuuf"���D;�w�}�ɜN������V�]I����+�D����47$z�e�򏜰ǐ"�_���ݡ(��l����K������=�&�� s}>�;j�;b�Ӳ��pf��c�rd����>�DЋ2���^g��j�O�Z�ok�<M"*/�����`��.z�5��[3���8�<ϴ����׌�a��a�:��;7u�5��MAH(�k��z:���:)��!=�	��f��&h2����k��q
O��k�v�8��7~ Ƙ����*Ɔ�r���c�PJ�a�W�Aa��EODe��<�
�!����YE�� ��Y �v���@#�6��ƃfZ�3��u����݋޳�����ԟ��N�٢ue2w���M�������!m�T����"�a��"�ꞡ��X`��<���܁�Yd���u���-������-��An���?4�Iv,�6Q2 G�k�:۳e	��)�� 	���~L�+�����P��^G&(���ń����v�Y⒭�m)4�n2��N``i����A����H��3)]k��NG���Xh�-
���#�+Bl�*94�P�1�p*��B.YR����4�K]���xS>uײ�]g%�dq N*���:eB����f}�!�N	��&Xݼ�3�\hj���$d��*��'l>>�> �/��M���;A�d4C�����m��mC�8��N��� n���^�tXt=N�qPt���ۉ����G1�,�n�Ds����ۡ��*<�K��?#���a|��[�/u��}%��9�3�����QF��͹������ٍu��3����Z3����H�O�����xw'?)`^���=1�֪R�3��fvZ���/�TA �_��o+��Y���ؗ~L�E�(���x���_eV�R�p�+��[e� ��j�t�H�H$�M	�ѡ��%�E�']� ]�[�˃��
ʜ<�K�����xp�=�2@>�Fjn��dl{o�o���щ:2o��/QM�#�����be�K��M�:��]����:��6÷��4!�~/���1R����cƔs��U"��q�	]-��6M�;K�H�u^�k�%�w�bp3�ZТ���4Q��8�G�u9Y \��fKI��ϊ(ٞ����PqQkC�ر���7&F�n$��h\aW7l�'�P�I1�Q����h��*n,�#Y
.��R�)�j*#�K�W��d¢�=��1�^��1��[���]����&����)��eb�<��f��m��j�9���)�Δ�.೚(Q��)ג���v��X�����s��?��l5�}��.�B��_��0�3�[D>hb׎[�Jl��~�(�Q��ζ�_���޵���%9�3B�b�d"`fn�~�໐�� �P42�$z`X_����*w�:�Y"�g�叹���~�����u�����"�Z��׿,�O%=�d���*�9k��R���6���B�AJp�*����a��aK={i3=L$�v�b�L�eύ�=���!�P�_IW'y\?����:����G�5�c:K�6u��j�7�1���#]o/B����ws���% �K{�/�\�T�}�ʜO#ʴ'�,&H�k��ڏ1vE�#�����uH#���]3:�h����b���0v��a�rJ������f֜�C糞c�7�D�Ɲ8��nIw_�	��V� ����Q6lͅ��{P�~Xw)2�wxI"WC[�	�H�ȴ&�Cj�:�G	`ks�b[0X��̛�!�MKn4b�=�}�^�z�K���2�RS]�R�L�c�D��rt���K�M\�Z�r�����/v�X���8$Ɂ�?�E�d�,��/]l/�PRdI+;Ъ�4Dʌ��j-�h� �J�⭻�]Ej�!�n��5N98��i�+�[��WDQT-�� Ր6��b�tL�ROJ�%���JF�	����s)�J915h�|���n�a�P���mB�و(T1)x=·�Obm��z���-���S�1J�#�:�=���=[�����Q^1&�����n�1S�W��byQJ��J](�L�L�������E2����,�Oi�b�C��ߋ&B��?�A� ]+�p<9EI�=K��E�5Е��o�d���xVP���2�����r���~ʆB�����u#cQ
j漄�<ҕ��J���ެ�~b�=Y�ޠ�8K���å
)��m:�em�C�[�a}�X:�������v?�v��5�=81%ngPr�_���X���(Ʀ��A+}���U.�U.�����>�m�u_w�TU.���|y?o�+kL��s�l�aT0on8�M�N���׳�7H�y������ �T��>���[y%�.�T�3r�;������Ԃ0ݴ�Ou�!U2Q��y ���ȾI���e�9	�I2�4s���.L���8N�]�fp�\	�T�y�\�	�jT�����/�ak��!�5dS�W; @��i�U_�̘8q��Ig��j�2��sR�ɛ2��/�������d����y�1qe��1����wc����r
�Ŏ΂	����綪;6��Nڙ-fF���f��c�OC<w3;���O��@��c��C��vF�Q��T�+Zj4泦W_���ՆI$�a��m-����h" �ԝ>$�#��D/���!EI/�5��%|�IS��Y��b��k�L聟E]"�ܠ���ٯ+���?3�uljє�W���
'�ރ��_���J�Y��a�-)6Ef��	�+T,�^� �l�"؝����z7B��K�i����)5�k�ε��{�J+�OKnCY@C�U�V $��]��.���(���E��I�urּ޶�����t�[���A4W�|�%!�"�:���M!	!� �]H��R�[��%�V�M�ɛM�Ɇ������ fZ(����&	���B۹����#� ���	˄~�
N�qҧ������FgԵ<8$��By�g�~����^$�x�A4�����<�k'\V�-�I�3T��,���d؞�j-a�ﯱ1F��³��Q�nM�]K9mrc-�}BT�޸d��n�u5�����bI�h�^J�"�5>��;�LCb����I�^U=��ٯ�c���-���y�1�{C ^ /t��;�䜡x��H�3N��p��G,G��,+�ѐ�ri
���qQݬ�F�b�����^$��0�\��;�=cކ��T5Ԣ�{/@�L!�8�a{y���[�s���dc��2��� o (�گ5'���~zy�Y�Es]忛�kXt���MԆ�8�gS9��U�\j�B�.4�i���h��?����ׇ�T0"b��e�o�4��%���l^�����=[�����y��<��Mz��o�c�����8�����[�y#�i?-�<Rx��չ�B�r����n��l�Ee�O��q7Z���7F�
�}q��*$Az�U�__;��0�-5���$����f�E���3���k��ڐ.�L$p5�C��gp�����>R�\(�	���>�f|�h�RႯɝx��{t�s1iؤ^C�����M��h��ƃٽ��萚(}yg-����w�v�W��e3RB;q�?ΐVM�/hL��"n�N�:��ƙ>ܶ���1�f#�x3e~;Aca���
]zcJ�ب
�/�{���:?�3S���$��|�tl�"�i���؍��f.k�ߵ6�%"D�!W)DRkS����G�բ�	ӷK/]ɷ\�Sq0��D�
����$��T���o(_K�8o�O�ģi�U$��k��s�@y�$,y���+�	���*�� �U��w�6]���a}W���i#�B.�<ȹ��X7�)CeX�Jqw���IѸX�V0R��ng��gcQ�<�I�QW!j�vh]s�N��8�*;ڬYÍ ��P}3�K< �@��.�\���:*�I���}�ד���T����5��!����*1� Jh�ቅ�68ע���h	E�Q�'�22�Nh���LvL�ь
�I�Y�����>yFn:��S����?4@�O\�5�����>\) H[�R�]����g����y�孧P�����փ	�u���W�g�r���>Y|���ߚG5.��A%�8"6_o<�^���W��K6�|�����bh�{���ԓNjwِ�6E���c�輫t� Xz�	[=��������	�z��*n�|7�1����lƳR��+_b�4S�M��O�c]͸� :)�}��G��{w��+�ﰠA�p�j`�f�mN��V��8�����j� �j8��Ժo��5P7F	g�b�'����tEq��w�c���q�!G�H8Z3��W�h3����Ͽa\g����8��i%���"�����?�*�U2����;����8B�X�8&(�0�������6�φk�;*'���@, �l���5��a�7v�n������B�"+!�)�uI$��F�]���p���^��yD��"�pޠ|��?�}D���̼��L\7r5���~�ꇃ�ߚ��Pp�쌫�Z�[|
n�bt�p�2G��W�q;c�a�ݦ�D����-������8���zt,��)E�Vg>F&I>>䅲��Gc!1�,�������8K/��l���F��PP�05q^�'n����U����g���>�n4���/� �����C�X��N�J��8z��H����U�k^�>��&p�㯫�ȁ�	ˍ��� !�3"oˊ��ܪ�	;g��	]��.��-%	m��6��v9�7��r����o�F�-�2޴�_S��;�C59�҄(�L �+���k"5*��@a;ݮW�3m��� ���@g-�����ꩃ[lR@Vd��rG*�4����P���B����zm�d����%��3�r
Fg�wAM�r�~h�4+z�u\�n���%��`�	[�9�5���7��&_�u��t�~�3J�l�X���X���JBYٟ̓���)�����[Kȉ�W��%7T��?����u��9��Z8`6��g �0z�b��k酸b1��o����*s���i!yA���������K�:{%�v]� J��2�d�q�3����J��:��J ����� �3�S���%h����au���t�\~���P��G7̩��� +�U��@�꫶��"`;M�5�O(��1 �j�w�~J�;&��y� �%�t|���ޘP*�WCAοV���8dB��W�#_�Lm�^��D�#�`�nn��ǰ�mZC�/0��>@�n��V���(��;���icx3+��)�d�d��4�Ӎr�Y���@$-��j����z����v�Yho�
Ð�x����v���0�>���۸3�I�t�MtX����4�멧{V�]��\D�e�_������6	�<G�(F���Cu�.��s�l��C̄(	����!�2L/Kl���[���r�	}u	�҆����<(���b2$�;Fl�}Ӓ!!�l�
:���G�7�A���� |P��%�Qh��@��0�i��l8�Z�(�a�u�����#m����S�����ZE��ߟs���cm��!�laU�t}��!�˪��}����� ���0��T\���'��df�v5����������b=4N��^ ��
z�=eۼh�^3���4C/U�n��f
Eԫ���Y�xױ�u&,�]� ٿ���o�`0�z
4p)����5�S����)*)&��E�mK���9�ʮ]��E���-ްP�5s[,`�����/B���mpOZE�a����dOL�'ɭ���F����+�;	
,��?����s��;��E�;�A-�ѼN��[���R����^ppy����^#�
�R�z.��۽X�p�7�l�Hh�{��îἚpi�\`�O�O�Tӂ%.��\��7	S� �O��("��%��P )H�U�e�ᡮ5���{��,S����MSk�L$C(��>��u�<=E]D7F��h3�1�4�i�J�q���`�}b0���2-)��W�����Ń������"�y"���T�M�z�[vMm�V!��]���c��`K<��w�����%4WNط>ӎr�a�"=�3%�냓L���
�P��l�ۉ$Q���-.k~g{4F��ڬ����-F��za����A� pZ����F�5=�Y��KquA�d�c5Ъ�2��)��$���Ĭ�UTM{�S��nmV#�斐��b�Z�C�ҕ�*B�c��wg �+J�̱f�_�ɦ�VDr������}AY]稜J�ԑ^�u�F�d�i~��Z�j��g�0�5���|og����I���rJ�h��>����^��s>L���Ғ/�sȁ/�xG�-��1M����D@�%��`�-�f��۲7x�ć���苲"^ 9��mg���Q�#w�R�� ����iL�U��;���-�+��� � ����M�(����:��=�S\
�Jժ1����(���WJ	!\��~��J*�c$(O�� ʑ�8'SJ���I�ىh���L���"�"�{vA%6����!s��,������=j#�@,p�fsɞ%�� p�-���`m�9�=�{`�#M�~�Y�I<�4���'{#0I��M�H�m|�:K����=�l���)�Q���b�e<l�Cʵ���~p����X�=��͆6D���ݲU���Q�?&`�̣^W��v㮘n��}��f���uE���ɂ��a��S��r"��7��n�d�<�S�?�_!�j��5n�+����L�J�s�y�lÃ�3�&)���=َ)����է��sm�j���o���ql�Q2h��w$���h?��,��嶏��#�?�5��m����xF���?���|�zJ��1ϵ� ���+
N� �q�����(�>�^UůG�N���V��Pv�L����>�i��|f~�mO��ǌ���t��R�bO���K�ԹL�bI�rK�M�'�z�����΂���]��N�J+#�N�,����=��Ĕ���&��(��WB󧺎���&sݓl���ު�p.W"��1
/��x�����,��%��#�5���SI�X�[���D&ó��� ��6I��q�X!���m��HǏe9 �(�
�.���e�`��q@緌�n8��'GR���m��سOü�����~ȯȗdJX�Y�:�t���=VB�kjr[~?X�wf�,������.�C����I;�d�9�8�1����-��؉5�
�Y����/�����/� �5�X�­�;I'#�y`�t������=�,���ږ�P����iH�D3		E!_�!�0dXo��$�KɄ��.��l3J�2�F4qn�o�{e�)#�r��?|�S�`e�9u����[�i��)6o��-.A�{""���S��9t���7~F:��;�y
x$f�&z��2*���Z��2s���ph�� r>M&��@����u�/�����15&���4=-{��2�I��o���s])�~��zv��etgP�k\���C�-�Bs��T��ul�2򵞿�r�ӿ��Ns��%�~�� ^�|�t�?��^aǺN�K"i}����7�Ld����{G�)����l���!�NFnm��k�~����y�>_H�����-Z)q Rr<�͐ML洁�H_��g�<��e:���g����9��`.Ē�s�����-*	�s@i�r]#������LB"-j�B>��)BzH��;��
�Y%��/�H�E�u4\[�(�,/#NE�������|����UI��y �����w��h:ھ�^#"�ǜ?6��S5��_O;7���~��)9j����|L��3�U߶����.���ݷIc��}���j�]5�'��B���}��~sp�ކ2��9���NE��l|��7
E�rw�	���W���Sc��L�⒯�q�'Cq';DW jw����vC@��<��E�K�(ET7�%ʽ�Գ^3S�/�8�6��+�/��c�9�M1+"�wzOc�1�Ǜ�`G�`�3�%�OyE��3�aJ�n5�w�'���U�,�29rx�i��|�B�;B�SR�~�ۃ�|��0N�_����J7�ʖ"b��d@����K��B�%f��ܟJ�A��̒W�Q�H$w(�M�%����"s����uj�f[̢=EM2�p��E�T��m��G�bAO��d�BU71���ӷ���n�OX?܄�I�j���.P��
��0<��(��G|� ��Y M��s4��Z�X� 8(�Z;�h�Bӗ.kK��p�>阓��Z���I����M��ŔAo��y�?
0}뤜�c(��������J(M4����KAME�����Pc�Z�������n9����8�<Vݰ1�D+�e�@��B_n�R��
�pn������P��EE!=���@ ���I}˕�Na�UAu�m�e�$]�����96�)g�>O��";�����&{	]SGte��^�(s)�������8�j����a���e�,)Z��Z�DT$X|�B�W�b�`��P���7��;��nFA��ԱdY�\��~v�ȽBVn����I��G��g�c���ߘ�s�L�Q �:H��]����x�He���-�W�d�9k�0��lk8�C/���!d �v��`؆W(Da��ZG��ˌ��s��!? �Q�*����g-�Z��nhP��,F%4��R���b	�t�6��!��ʀ�_���i����\aHiU��[�=-��c�~� ���tc�J-�v�<�����
r텾�Y�;��^�Q��_f7�f�;��bdq��:�%���se�Q��sb(��Aa)N� mʧ/j-`ˠ��K7�zY����~��.�!I��L0�5��k)!�/��Z��s!��g3-�Gտcap�*)�W������M*�8D+^v?���B�Țuy[U�]Ɓ=o"�����|x�Ah���E2y���J��.����䎶;��?(Hu�1�RGr`��B��~y�@�l��s"��/�:q�|v�5h����$w�:nn8 |p�wVF٤��d�旑��AEݤ&a��	74ےO,$9��ܼ/� �8�G�Uu[rI��L�+�/�E��N�<Z'�c0�tpo���4����Q�g�
�#
�nZ���]�t����)�v������h^Q�A����;�i���x���o� iq�um�����JݷK��ں
y����I��k���}O��jK�3��4�)�I�Y]#-�
`���I��O�C�T|՗!_��'/�%4�eր&�n�� @m�1�P��N_[��9a�C<ٲ�\��9ڄn?]�;�!�䔴� v���f(���!�do��W�k�c��%��+�~H��3��>�Y~� x��;��D���:�N��J��}�憒0/�E>R�X����w�"�i�<�vk��2�n��j~����x l�t��l<t`4156ы��\�.��Gcw�f��3M0��u�m�u>6���:���))��T���c�B1u��@u�\�����瞒��އ�3 ���6��-h��V�e�ӂ�Á����Z"�����-D� @VŇX���ߎ�`��_]�4��BMcLAw����XP��2i�X �^�Ehc<B>�l�:�1��\pЀ�-K�a�����g@��bB�p��1� 9�s=Lorߘ� ���Ҭ��|Ot�)p>��.�4RO���������@�&���T�P�(����S�Z�<Pj;��^����6L<���vg�`Bz�8R�7�?��V�����]��]���BŦ4�F�e+��νDF��Іϰts��h��(��l#yNH�Nc�.�#=R���_�S�0ۭ}�3�|v}V/l��K������&aXy�N�u��G6������S��t\��d*8���%@f�~y��AՈ�pZx3*�����e�l,����|v ʠ5.�]�Mqd�O���L�]C�sdZ��Y|!�Τ�<w��ir8��Aj��� 2�c�Nj�Q�;f�9�N�RW	|/�T%�bAD�e`>XJ�x�Bv캢����М'
�.�X6s����b��\/�`�M��ͣ4�F��-9�'��0��|)&��8�����vf�P=W�>�ҭ�f�wчRA5�dM��ٸ�|���J,Z͇���a�Z�y�l�U�#�1$D����r��an���X�>ʝ�]����_|����=j�vR5��Avj�e�}O�jd���K��uk���ҍ~H��`��#Y�\�S�)��[�+��E�,f�����P�l�6�9qp���"h3��Ki?qu�ސ���+��=Be�PR�� �Y���#@]Y�c���=M���ti�[�f+�CT_lF���3�f�Y��X��8W����W�7�]�N��������������:�jE�O[�f��e�y}� �}�o�a��y^�;M�f1;���r^��NOK�o��=O��&�(҅i~\�&��z��(2��w�t�J����]էKO1�K�뽑�}z��3w����\���pO�!����Ӕ��ij�\���EW1�{�� �3�ǜ|�Iձ��&���(K���3�5�-�Č8�Rt$c;��4jmT�Ɓ�)v|��/� ��l�K��*���������ڽsy�ԋ�.��<�`[�l#8򧔧�ѡ�]��\�{�6��~	�|�X�ϑ�'�<2"����c���WL�H�=����a��X�GRm�Ai�[�5'�O�ih���������]ۭ��g���?�-�<~j#�S%�쟉�MC���3�ɦ�ٟ���3��v�T���{��Q�6Hd �&�$I�xb�ؕA��,�m��Z24�f�Q���q��!���i�Q	���%�TI�X��,&e(.��6
�VXܕ��z�*����@{�E���g~�c�'��Ji��XBSvLڹ��B�m���a^A�N�y��`�3|���3\����K3O)�k�N�*4�Mi�/, |���Cs��a����bA!�Ot���;D̠��_�>�	��-���I�T���������y��	��"_�o��p1�u.\n{��E��n��3�ؾ�ȱ�-Sqlj_�]�mގ�k���r���v��<���W΍�U�R���\C���jo��-��=����+��)-4�/G^q���>�q��?���Տe١�B���	(��