��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�w�tܔ��@��zATe\��5Â02�}���iL�t�F��������T�NY��y��ti9) j'�A�&e�U( p���9��C�z)N�`�+Q|�w��i��Q̍%�i$NzUC�ﾕ�z��v�K,g�%�zI�_��j�\��u�Ǩ��.�}����	N$9|���%פn�#X�1���c�3�����.���V�e��-�lZl��c�_`�Ƒ��#�R5,0�0�VǓ)
R�Hh�IС�!r�0l"��g�joyi���ΉY��1�/^}�E�s�(�w�fW���8XF��vC�v����\�e��&�>?P4�~.8��./��<0�9|�`e"�kq��fy�� FƗ��ے#�7ٙ�=˘HCф�ڧ�$%��eͨ���~wFfLJ��m8��΀���dj]����2l{T(S�`S,�+؄�VPye�Q_{��?���3���ӳ� �KٖD2�a��|������`=��I%�nAD�i
��̝���z���?���2_`�#�7{MU$d�a�4���5��vn����#��&i�f�B6y�J��y �`�n+� �(�!?��q���$޹���+�;��m!;��R��������!���$�����i37�$GX���^9��n�x e�L��l��z��S1ڢ�?�/6Y��`��f7z
�2���;�j2�ħ�b�4��4Y��=��k?�!�sQ�h:�((��T^���@��7���8�Cyzby@��-����t����Jk���w��­���<�,nmT�R ���>��/`H���"lݺ���UÎzP��!)']ޗ]bz�/!�̃cľ=X��sg[+1;��ᯧ�s!5��U�x���/<SYoU.�O��&����O��.�vu�ڑ9�*	M�X�z��-����x��#a��tY%���6�Dc=?>{�����s ��,2��X����3��d��F>���p��F�ᘽӂ�é�j�2�Y�1]�5��
g[B�B�p`���� mq�_�~��y���C)1N
n�mB ��'��[!�����m̘�������	`',!��#iyd�yB�^�Af�ga��u���Cdjm/����T�c��G��s�����A=��YȰ6)� ��L�jڻ=��d-���|/�4w��!&���<���Z������[Sj�̤�?�[��	!���m*T�S�C��z7WGvYܕ�΍Ý�`��i�|�
o&5 ��z��7��{NW�M0�z���}1U�FF�|�(�Rj͂��2ss�����Şg�m�ݤ�^�W��ږ���e�����=��� �M�H����F5YS�]��wh
���A0\RG2k��d|d��?�N);���W��	��Ɂ�s�r���}�)1*���Pg�Uw��oJ�6D��L�H�f	e�^[!`>X��e�6ƽ�����$�s���q�9�Y�Û�L��<�3����o�[� :]1�U���q�#i> �e~s3� v��Ä��TB_Ż�#��D�$	3�i����	b�x>�Ǖ?_��Mͮ�PK���ZQ��LF;5� |��/i��v��O�1��5o�ZX�