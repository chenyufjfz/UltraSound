library verilog;
use verilog.vl_types.all;
entity controller is
    generic(
        SIMULATION      : integer := 0;
        AW              : integer := 10;
        DAC_CHANNEL     : integer := 3;
        dac_pcmaw       : integer := 10;
        COMMAND_PACKET_TYPE: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1)
    );
    port(
        clk             : in     vl_logic;
        clk_2           : in     vl_logic;
        rst             : in     vl_logic;
        trigger_exec    : in     vl_logic;
        ctrl_in_udp_hdr_valid: in     vl_logic;
        ctrl_in_udp_hdr_ready: out    vl_logic;
        ctrl_in_ip_fragment_offset: in     vl_logic_vector(12 downto 0);
        ctrl_in_ip_source_ip: in     vl_logic_vector(31 downto 0);
        ctrl_in_ip_dest_ip: in     vl_logic_vector(31 downto 0);
        ctrl_in_udp_source_port: in     vl_logic_vector(15 downto 0);
        ctrl_in_udp_dest_port: in     vl_logic_vector(15 downto 0);
        ctrl_in_udp_length: in     vl_logic_vector(15 downto 0);
        ctrl_in_udp_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        ctrl_in_udp_payload_axis_tvalid: in     vl_logic;
        ctrl_in_udp_payload_axis_tready: out    vl_logic;
        ctrl_in_udp_payload_axis_tlast: in     vl_logic;
        ctrl_in_udp_err : in     vl_logic;
        ctrl_out_udp_hdr_valid: out    vl_logic;
        ctrl_out_udp_hdr_ready: in     vl_logic;
        ctrl_out_ip_dest_ip: out    vl_logic_vector(31 downto 0);
        ctrl_out_udp_source_port: out    vl_logic_vector(15 downto 0);
        ctrl_out_udp_dest_port: out    vl_logic_vector(15 downto 0);
        ctrl_out_udp_length: out    vl_logic_vector(15 downto 0);
        ctrl_out_udp_payload_axis_tdata: out    vl_logic_vector(7 downto 0);
        ctrl_out_udp_payload_axis_tvalid: out    vl_logic;
        ctrl_out_udp_payload_axis_tready: in     vl_logic;
        ctrl_out_udp_payload_axis_tlast: out    vl_logic;
        local_ip        : in     vl_logic_vector(31 downto 0);
        pcm_udp_tx_left : in     vl_logic_vector(23 downto 0);
        pcm_udp_tx_start: out    vl_logic;
        pcm_udp_tx_total: out    vl_logic_vector(23 downto 0);
        pcm_udp_tx_th   : out    vl_logic_vector(7 downto 0);
        pcm_udp_channel_choose: out    vl_logic_vector(7 downto 0);
        pcm_udp_capture_sep: out    vl_logic_vector(7 downto 0);
        pcm_udp_remote_ip: out    vl_logic_vector(31 downto 0);
        pcm_udp_remote_port: out    vl_logic_vector(15 downto 0);
        pcm_udp_source_port: out    vl_logic_vector(15 downto 0);
        dac_signal_len  : out    vl_logic_vector;
        dac_cic_rate    : out    vl_logic_vector;
        dac_run         : out    vl_logic;
        reg_addr        : out    vl_logic_vector(28 downto 0);
        reg_writedata   : out    vl_logic_vector(31 downto 0);
        reg_rd_udp_mac  : out    vl_logic;
        reg_wr_udp_mac  : out    vl_logic;
        reg_rd_dac      : out    vl_logic;
        reg_wr_dac      : out    vl_logic;
        reg_ready_udp_mac: in     vl_logic;
        reg_ready_dac   : in     vl_logic;
        reg_readdata_udp_mac: in     vl_logic_vector(31 downto 0);
        reg_readdata_dac: in     vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SIMULATION : constant is 1;
    attribute mti_svvh_generic_type of AW : constant is 1;
    attribute mti_svvh_generic_type of DAC_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of dac_pcmaw : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_PACKET_TYPE : constant is 1;
end controller;
