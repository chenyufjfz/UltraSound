��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>���q�;�;�g�?�_�q�-�m��5ʞ�œT����
��cFZ��R:�'��o�xE[�I�N���B0ˀ�2|:{4�C[�p6~��n�?�Ϳ����^:٘�!,�i�dF��<<���0������� �Z�=+C�r�.3]r�p0��ũ��׏E�L]�kvB'�w���f
c9�v�F�=�$бK-�(��/s7�jج���l��'s��2���[�=H���O�xdP�=�|@O1pJK�~	0�='�F�;.7c"�c�DΣ��t�{��{t��Vœh&���ڝt���3�� ��8Fko�@��G�冕L�!zx %l1c�l�^��$2�;��I��}#tJ�I2G
��e�ό�_k.���T�p�#�Z��(n{e։&�Wd���l� GT� �"1j��y�yT�!9��-�*����U�vi�e�;U����EyT;��ª���S/���{nv��P���ҍ����S�-�^US�Gմ��������@�e�ۉ8ݻ]�]>��(�����F�q��QF.oF�/ �8N�$5�i3���&����K������<������'�An����q{�Q\W�?��zb�Ӂ�&���4GJ�z87N
� X�X���@��"�� ��͡OmgBBk�c��E����TN-6^���	���+i�'ֽkYnj)�� ҿ Ő�����=�鶱�5yU����5��2pS)�r�n�ߕXK�wj_�h�U3yun��+�Q<5�OTI�Gr~���-'B׎��I�p�})��M$�,fz�ڬK$8?���\�+�� �Z�diDkJ=N
t���E���rD �9���d�1���+~��G��֓m��,��xv~���x�J\E�b�}Z�����Ҽ*k��
2�����wѮ볜�[���Gfvք��Dڦ�;�Mq����z��"��4:����x��s?��,#�E���¥�q%���?f�
IIq����p�"sI!�8=�}KN�F�}�?U�&�^ʴ�ĕ�8�#�R�(1�����Xމ��}[K���I��M9�!y_E�_�b�ś{����n|�9�I��R���مX��<Y�ޘ�T��B`0�M<ţ���Gj���	�F� |܇|lʚ����ܚ�R���AВ�=�b��0�n�_]pTw1�t×0�4�Ό����s���z�Έ%����I�Z�>�^�m)���e�U<ժ6w����
E�*������`On�9��&{<4k�u�w*��V��t��2�Uw�B�[&�K3�=O�h��6|��-l�VT��b�|W���/��t���Q����t�T��9a�i�(\���x��_�;n۹�ig|�<!�����+�w#bi��O�[X����C!�<�J�����2jng��@�la��3 �z5��E�;�k��n�7�*��
�A���4X��I�v�B�s�e�����p��%e�p쵺M%��p�a8fN��Rk��W~�����i_����U��9�kS�~m��u�B��o`��6O�}�AI
�r��'����=B���pX�5d~Q�-i�VsY���r�s��B"��{7e&B˲2�m�o����F�Ǉ�.Ɋʗr�;\�D�^���� ������.wP-eq��Zl�5�I{��ϜA%�q�-\0gR�c��6[!�����F�|HՕU����o\3 \N^��C�Xm5`&H\>n0��Y$��*�9ƣ��G	4�8V����`��Gv'�����枔�Ab'�������f;��91L��I��c,SS(�zp�#vĶ���C��@��	�/�g�mJ��p>櫄Q�e*�Y߯�{Ǩ�ҟb�jח��k��0;�ᒴ}���ġӈ���EV��5���dA�]Bu	_^�B�A�i�a���g^�uW����xF\��ƅs�y�2m���,��ՙ��tF}ۛ���sH�4ʱW��A�m;N��;}�tY�r0�����.F�C��#��":�alvbp��&��?͓���D��~��J/Լ�y�@{�UzݙH��_��Q`�O#�/̞���~�y��4����f�|��-�4�������ͩì�7�;T���`�ˠ��Q����-��0��H�{D��D� k](u�����3	F�q�����QSg���>���iE����<�,PG������|SJ��L�6�i*{��.��l�2����6 �K���7�G�����f6��O� 6�++�N��*f<	.y�d`S�Q�G� $�r�L���
g����\w�OJ��� ͤ ���t��<�9��T�~����KE͸�`�鷺�!�$���?�V�5�z�˦=�ܣL��pk�c!R�:�}]�H�� �'��BB{$��^̠�=a�VӺ��}�hH�t-V�ķk���O��'��DB1l��\�^���<Ly*�g�cNs��FQr�|��>^�������&%qIW�wn{ы�8���򩿘��Rj�ƽ��
%|e�y
k2A��|=k�Ȥ䂔�B6�[	�xxiVɃ�$��J�p�����ȝhÓ��"|Ӎ-����.��|�����h��R�Ӂ�-Ҏ<eᇚV�`��]e]�<t�ԯHl�����E������A5����H>"8�_�5�ze��*8�8�+
�k���K_��O}V8���[�v�{KC:C�Y9�H��؀�!�9̠�QS�J*4VWuc4Q�щ���n��u�ŧb[��֛F`D�������!�ج$�����A\`�s/y7,��S/4��I+e��p֪S%o\B0��=�)�5yA*���������&��U�Z�Eu�l�T!���П����̀�gc���L�揨�q��ǲ���i|9)�������4R�(��W:�i���Q��E#�|%e�%�5�����zeP�A��ȗ|��{��F��W.̌2vl�6����q-��i0s@�Ubo�P�/�2�F+���$@�^����TH�HЬh2���C����}�2o:�j�
��_~�x81���ˍzl?���X�ڱ3�C�t%{�ؓ��!v�}?O��`����?�:j�Ԟ�Ԅ��
�*�5��V�i�rdM!���<����p.T_�mt�`t��ոwSz��ŷ���z�B�".����X>l`��C,u���-�DW,2���3s_t�fe@y j�`�ɩ]x�k(v������e�^'�(��Y�[ ��р=����\���g���c t����}����ZF%��ƔeMs�Y�*�ȩV�u l���¤�$��ᗟ1��X�:��o����j ��7?11�D���`Pt�o[��\�\B$۲� ����p���8$7�~�3�G����]̂�N|H�*��K���K�?���@ߔމ�=�Wa����И[�>�sZ	�9�A��,!ND�?�6[u|˨�3ȉ�%e���9����C	�Z��,��O�7v����Q��w�S�R����)�����<���5K�!�po�\��!T5n���݌��2�n�� ��0'�V���*+���qQ��H��W��`�	cb+a��I��~���_���^�C�J��w���0 �FSYV�&	�{����f)��m��R&��}�d�jP�g����L#�o(;X �������Gn��e���k�:��1�_>M+}Gk]�Y%(��	�էf@�	}q�,-�1~��0�\�?��	7�o�������R�;�l���Y�/�w�G�����	|
���� �Uu���������	V���5F¤k�tTk��;�@�!Ņ{�Ä��E��r��_
����xD5�&V�M��	^��C��!�Hr,x�Z��6�:uN�P�99n�w�\����Zu��T�c/2�Gn?M=xy�|�v�A�߸�
����YJcDO]��I���S��0�E"n�0M�=���|5T;�������<���5?��Ɯ��@\wk������P<�l�}�P�]��+=F� ��'�E+�	 d���ZFw�=)Ә��W��:[$Q;�=��/Z�ue�P���hn�K���}(�"-���9ux���ä�:&Ӵ��e��e{�I�ݕy�ɳ�-Rν&>��NE���m�
�?�GH�W�E'�ۆ-%_����G�8toc�@	;��km�M�`�m��X�c�7�'�8�
�sa��O�2�rh�0)�*,�F�p���>�c1�}β[z��nf �M/얜CW��q��d�m,����G>5�Ƌ����I�M�k��N`�5���W|�D�{��[�v����	����.� h�ޖz,������E�
�i�� �"6�azU'zb�w�Pɂ��8�s�����3�r���+k]�[D0�x��Ї�e�=���V>��<�Rf}k���J��A�q�i�G͋h.�I�!��{�p���䜛��A�V���Z���
��Ҫ� �F�Jkس1�%� RR�[��j6�M=Ke�\F����*�M9{4L�&����i���*��s�MA����� �6��̠�� �'c�2xME�����HFC�cQ�X�R���w��t�<�us?w�}��L�r�O(���oF�� �B,�X7��d�|g�L�;y��q"@�Ѽ�,�u�`P��]W����F>�V}8i��k
���g~l
�Ď�>��H��Չ�������������CX�y��7%u�|�m�����zY��N����mb0.�B�y|��s�h�-X������2��R`���[A /=E�ߚY�YIv}��s�c&��>����#�۵����P��U�ڛ�9ׂw�Qyz��;�E��ζ���c����YQNF�;��"�I�r�������z�%O'�Iw"u64��vg�����n�ge��]d	8vaIν�Ǽz����c����:�]z��*�~�q�е�,�!���t;$5�iZ��������|H�и�
zJ�<\�� �Cڔ:Hѿ X��_6F$ש�~Z���8�h������J����ϲ#H{H��ġ�y�GB22T��2h�úf������Hz	S�L%m	�SM�ߨ��A���8��id �p�� 3M���ͻ}�z��X���������Z\��;t�|���9���?'bN�Y�-b0j$���>)��&N���}Ǚ\m�L3�L>~.#���^�������#(w�d�{6( � 2#Iתnڰ ����OպI �P��\q�R	��B��H��kz�A5�=���Y�I���n}��Tu���
9���/Ln��z�t�HR�����L��4c���u��;>���R�!.���'��4�uՔ�m8RwΦ�gg�������j�n�֩~
��Mv�ncP?�s�_l�:�e㻼��z"!��:~0����\\/ů����~ ��7�T`_)FH���S�4~qI�����z��:�����4]#`vnh��{�(�J�y�ǮO���Tɻ�6�wVa79O��T.}؛�SO�>}�p�^y��
L7����rS<��xE;&A�~(y��D5	LB��b)V�
[��
x�K�WW�"f�촺)�N!�S��gC�ᤕу�bR�U�������F0���o\Ɛ�H<�˾�0����R<k�����D�eH]�Z���Wt4d�ǰS�`*oo��`6Y9M鷒,�}�����n���`��'l�	��������ֿ�,�����L09����@(���&{L�@��Q��y�l��-zj���U���4��׹)���������[��Y�`�F�{OO*�m��/	����S��^I6�G8�� x�䮚�7 C�7����~�qb"0\��a"u9A8�w��+������Ϫ�`Ӕ��T�j�Ҍ������Z�QѸvq��3N��c����c�X~wPV�aBhY��3�kߗ�)`�g���������Jm&�Qh������c�wX&��|w<b`��[]�Ä���T�2�Y�b��ۆo��i�C�G����$���R�~�!��&]�s#�,�T����?[�a0O�L�r(@9 �Q��j?lL#�Jl�d��ə��Z�E
w�Ev{#7�Wٰ�y�	ߕs"[�p��ND>Wy�n3wx ���i�	̸t�do��`Ÿ\�EϮOU��Ci��t�"���q T�� �Wp��l� ����;%��y���&��&��75���j�r�#p��b��;�Ϩ���-�^{���W����G��1�$ll���}���Er
�0��C��z����+�F�9_p붑���'.N�,��b�sF6b5�P5-h��k��~z�	�w;4r�ܺ��dg=&_�ٲc~�SX�t��h3��I.��+S�Ҧ���h��c���5qvҷ(�5�n�=���UȲI'�Ӆ�[�/��j��X�|�:?������m�6n�eu��;����>`vy�����m����2�ExL����0^"�S��^����PO1� �_UM��������r���o����}{�/�\�,�݊�dC3c|���~��	B�9Y��$e4�$���v
����1c�7�Cy8�L:M	\����9$��)��6����S)��k!�!
T�50��l��La�����o��K!"�.O2q�ӣ7!�Z�'�:N-��S��z�e :)�Q���z�>�KM��J��c�0��W<���J��->�̦�q���������*�É�ɂ�oN�i4��F�˒�In]X0�m�W���`�
l� <-E�ʓ���!�ՖS�����&�+����ï�\p@�iع�ӝQb�U��3���p��t�t��O?�#"P��/�A�G�S��8��D�g����A˲���NZS�}���^z\�����>����U*���"�O�@��[�����Zs{�:�GN&���ƱU�;���ӊ�l��F�VB���B�X¡j�j�)@o;�P���S�Th6�)~��=���!']2XD�'��s/����Z���+�Ӭ�p� �4o�����l��.ΗZ6��	����{�ñ��ݘm�AsƐT��q�6"�(���I)��9����h�ǋJ?�����%��/U����	T[��ݔ*0��5B���Xh�/lg?q�D�m�L2�	����P#;�("l� �AX�Y=xuL%1���Q�K̈́}mꈑ�<o��<nJS�0�j��F�8ֵ��v�����G�F��V��<�F�� z�r6�������F�y�I�(� ڕl�+�r��s��OX��f���^�.�.Ӷ�s��m��0������!@N��A+�[��N@U�G#Ub�
Tv���?�/-�t�Ւ5���W���@5LC��X�z[ r$QNI��P���(��e.�ʰ�@B�?�x �k�'���_@'n ;�Vt�E�?f6�q	:i���E�1-2�V";�i���J0���b_��X�!(����j%r�\?	���z�om㦈}�w��ߛ7G���qJ �����a����u���������`���f>�9���>nL;�k��aI&���,3Ir�y ����x|���� ��� d-E6!�Q�;��	�%��Һ�`^"C�+#��!>�?��"ɠ�:nؼ���R�3a��Mݶ�9#��p�+$���sJ�{���y�b�(��o��*1�G�BhF^����j۵+����s(��t���~K��{H]��P�Z��T`�P^$����a�o
YY�W��
��*(zQ�� ,	:=V�Se{��x'��������
�O��U�<��Ua�i�'k�[B.O��q�P|���Vz?wV��h��!8��ADY�lUsP�n9��S|���4��T�~xÊ��ĝ{~�J�sщV��zcl�R�7L�c��
��B����?zƁ�^�G�b^�gA[~�8M���b=���M�B�v\p8c�1�6��P�.
�@h�W�]_Cght�O�3<Z�JPQf٥�\ ��~BH�E�-�R���?�;C+�d�J/�C���~�e�2X�?�c8�hP	~6k���슩��_ź����c�f���^R+����b�(Pt��_����PPz�d?�tH>��lQS����!�$-��BD<��qR�n�ɨ�f���3��a� ���a�+���U@�u	�T����\�B#�D&���AK� ���}wf���^�ʕ@�+uc�w;=�Z �]I��@Z�E�� �ܹu7��ja�ț� ��~��jB�w9�����F/�5ir�`õeSΒ�4H/�٘Ս�&�s�P��C&�"����9�����ad��� h��3���Ra~�{n�B�g
:�G��[<RO7l��,�����U���I��ߥ�%�=v��ltkz`+���Q��A�V��@9���\����?��Pݥã���ؽY��W�G��Z4���*t��*W?M�V\�J\
�S�%:CI!��%:^O���n���L�|y�,EM��_�	C�S�">�y��fە� Y��졦Rsx�õ~'*��Cd [ޤ��庩���CQv�`5L;��Ṍ27`�\�C�'-�9����f�1��\�j�k(Z�t/�E�>og����W%� *H�H,�%�:�V?�����׋��@Gk3���uB��Н�,�)������M�W�C�WK���|�_y�_�i�{�J����ә��+�g�'^RtO� �����[�&�0����ƾ�N�F>�f�R#ˍ��^��
��3!����t�)��{h�}b}�?ՍT� ����l�j��X�7�嵛f��y.f��o�OZRCq��>(�)΁��~���0�{�k�gF�P�����u��������d�|�|���ף~4�����^��� ��7�L�RV�ʳ"�➮Y���Q��*@�dB&�ݾ��"���	�*ͷ�   ��5̑�PZ""Ś�!�����۽��(�g�͛�
ļ+z����+�w����-';�f2�Od��$1��G\�܇W�|��E?y&��ai��j���X��7��b�oܔ tO�[?x;�m�d|�Rf5Q<����r�T���7H".O�)^��'l��ջ�m�*�_��a��rq�noZ���#�F8��j�����H����FM{�x�A�fV{:iH����OP�sz}7�N�GM���|�b�k�ZyⰆ:ҹ��4ƕ�!��QeQ�:�1x���}b�������v1/���x
�HlƹwQ��H�����g|�	�w;&��1*����()�7�̺=�GNt`�g[�>�,��G����7���(9�]6���~�a�(�y `1�2��~v_S5��+�nP�>q�Ը�D�<���&��x�j��JSk�,r*L�'G\U��K��t�s��a�����q3�u�%�4��vR�[UOҐ��SEk�K�߂k���
��	*�2#MVq������ėƨ��9��%]��*,��1!^�,�5�;Tz�3��NW{�6Q�'H��>���M�V#��#->���~�� ҩ��cyڑ�N�~�u���柲�������M'ѲI� �~҆�kh�����c�O3���,C�@+�̄}��C�� "je��8~�R���>��=N��ؼ�.nT���/�:��䣁y�~,�{��?�����JR�^�${�@�_M@�^h��������kL��eb��5�t1���^�hu��=�8WV1Ȋ/b�I�ϟO��@���e9'C�����N�#�ȠE�A�53=4hf���};^*d �a^|��c�B�h�[��2)
b�̃�>#4T�&��K���JR��_n&��C�+�P�B�;���MT	�.�'���)i��B��d�:Պ�C���+_�tV	7�N���gJŵ{+�$��?�r��UD.�o�S��v��%�/�Dp�{k�d�U^�@<�=�r"�Ԗ�[�h�H� ��$��Щ�ت(�L����F�b�M<��3����慺$��������En�dc��m�^��-|�o�P%�1W�LJ�[~�����w��R�n�(ט<��"C��dt}���8��X��*_�_�ۚ���?�0��K�n'��4`��z����`W��W/��@�v k�MF�w�P��kA���Ά;_R��9k�����i��z���<ՊGQ��T+��� �Q1"�I�ze����@m	�w����uO�ō]�W��G��r�`U~ފ��mq+YO|A�;e�-)����[w�쫵�h�s7r���;����R�Χ�NͫX4�RYB)�y��c�K7'�A���ӄ:���#b|(&G��IP�c�a���&���Ž�>��a�~[�`P�%9�e�
�sU1 D�/�p䮄3u�w
������w�8�Uj���Իٙc��c+���U2���w!'�d�2��i����LjS��]8�Q��8^����J%�5P32m�ꗴ����������E�#�$"$#�řB��˅ui.�k��\.�����PI� )�11ׁ��FN���Pq���Q��)����HadQ���Dh��Ub�gck~�|tb�����g��(~���4�|��Qe���c.�S%9Kg@]{���(B����:Q�jFn�ܤo��z���b�DW�R6CI�����ھ&p[1CB(�׃���:#j�u0>�G�h� I�
���I�EB&�ɂy�\<�Ф�}U�����mA%��!'[8Yɠ/5I��c����v0��3mЉ#�fLs�����D�fKˊ��)r��MC7:'�AM�D3�:M���� ���"���yfyD��B���e�P���LT�	+����X|��RcC��x�^^OcO��8?���r��ǈ�S�+u�JX#-z˲:31�{���Օ_&F����v7�2i�[�k�n�J�kp539�6��xxfo�	��������0v��8�rS��[�
����KN,�z��r#�������+ր*��L�6����zjTE��1{���o œ��|%��F���#p:"4�����
3���C��arm*�3s�$�vʾl��K1+pϪ���Q��*\'��.��ٷW�E�9Q��	n,>�5Eq8/?���Y�켿{�o�V���Pit�4t���|'�Gko��5liD�&(��L,s�Ͱ{���'�UUB���Hd��Ib���~��J%�8���OdZ��ٽHI�zoVҖx�k���]�VtѨ񟊥��W�A��=��������J�����_&E�@l�-`|�Y�%��pu�[G��2#�q���.Ğ�2j4��kxCej��$հ�qa��$��hm�"�����3�`���3}�G{�G�sդ�-p��=VB����h��o��M�W[!�pE�}��|�ni�dC-��:�f'�m�����ŏ���p���N�+;-�0��~�F�~��MSV}�s;O 7g�� �
�X�H�|�|.���_�2J�fX%���8@����Q�q*
�n�����>M�`D�x��D���lT��dY`�@3Գ�Z�d������Ru��Q3G��Ϲ�BU�����A7ǲP�ĈEԳ�
��	�zA{u?n;*kT��~LB�!����c6�Ik��? ��e�����*�=RFtX���h�)�@��@�|v�Y��KX�GG��-��i|�kwC�2�����I�N=|�R�g�����LI�Ȣ�`��%�Q6!�_�ߓ�T�Z���2�����`��>;�������K��/�Q*�G{�&W
���W{ |���ͶQ3�\��Fꆷd����E��Ɨ���p��w�	�s�Q��E���z�kn�`t6�$�IKF�:�;��Z�\4���VC�Z�Laֶk
���Q�V�bk�� -=F�|D&�,��*���Z�Ԫ�y
%N�� ۖ3�� �"J�8@B�By�'��(���c��b�lL�ވ���oo���(�!���v��o��{����Y�J�"@!!?}7�[N�aN �ܝ{ǣ���@�[B�b�}��H[uw��5y����4Ok��J�B�ǚ�'��/*Od���y��l��c����
�u�I��|y����{Ա��^��,���~���`X�8�J��
K�v`K�[�s�H���=&�;��c�eekP?O�K��_�V|\��ӕ,/�6@���7��k�P,�̻D/��<�9Щ>G��Kx{���`@V�E�������Z��3)/Fϧ8{X�˿���˚U>�Ű�k�v��a�J���&�GܦOA1S�~	k�M��"�����T�w(�7_���O��2WBt�'e�y`�@m�=ٴ�s��\$/K��{-q�߶��z�|8�)aؓ�4��d��/�.��$tx� 5��� ==�uQ�K��G�����5�t� #x�p6d! ���qM=�L��ʌG=
G��{r�&����Ĩ��頡?B�{���#/�$�����uR����uj��7���#Y��c��������=�1Y-8���<M�N��<d�����ϸ�U�R��J�qφ��s�ke.0�i��Z�0�k%�UM���13}� �%�SC���
%b�(�0�Wsjp���hODJ��E�L�b�]�S��Gڇ
�@�UWz5��-a�w�'�w�*�~�bB}��U����?�2�hF���}I>͟N�v�}������5�G�֔-��+a��/S��2u�Ϧ���4�Ŝ=g�ǹg�c\Hi'�#�lQ��;�f���/d2�����vRX4Z�[��� go�o���t���J�|�ؗ�q�3��\i\o�ȉY�B� ��R�����C����yh�n_���u�>]Ek