��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv t1������O٘?�)/;���;�+	��۳�c.�Tw�R�.���js�w W_�k����|���vY>j<R��ZL�����X�T��ã2�ސ��]4x�{
r:����_z��F��Qq��uZb�sG�rv�Q2����=�Ђ��&�=�J��0���������4#)2�}���mc	�NhAk?nt���'|�3��bTJ���+�~��E��{�ɷ��)kLD� љO��?���2�n�
W�ѥy��}.V�ߡ6�^G�&��m4�jL��e9���M����O�7�js��!vf��uR��k�1�+����\�m
�.\П�g@�� �ET�"-W��A�4Q�A:~��e3XLj�X�buQ�!�ý�i<UC$d�KLW=�p*��-����Xw&$x��`�"�j�a�}�n���H�K`�B7{/�{0��k�ͷ�Ȯt~�$jc�)f���h�O˄\��p�M�kܒ}�O@?|�P�S^�m$�|��C
":�?
2���~#J&?��6�qi�z3��,�UT��F�~�t�N�%)[��#�葚N�ъ
�{��aJ/����Ѕ�f�z�7
G/� �3���q���9	\_QB�t��Tp���Y�Qo��3Ĳ�-M1��Ȋj���}G��7}FS�R|:FK��ͻ�*\cRB�)�H��7wt��ü}��9�Wn��W��ŗ������Z�����̶�&Us�c�Z��q�%���q&S�n�[&�fP��x1G{�b��+�t��+Eq�����6�Su��Ru>��a���Q��[
�0�س����[�;�����Ѩ�&�$
b:�ی&�j�$"N�$vp�"ݥH�lo*�RSE�+h���Ʈ������,�����\��ɣ���xwB.�̑�'U�ѥ���75p�����х��D�b��`nDa����E��J�@M�X��E����P1� 5�[;c��a��f^b�2B�E����~h��<�C%����5Tskᔏ9[�����)Z	]Yfo�I�.Ut����Жf��$��$�����F�(u�,� uU�U�`/V�fF&P>��_�C��6U�>��M�.U�����:�eF,ʏ�D��m�3�|��n%�=pC�b���M�	���U��^4����
��#r�w-�P����&�K�y=<�8�ք�������AY�mX�6���3�
`�}B;�£k��Y�'�Au������Hy4 K7�]��?�?��e>�5Ђ�mX/r����6����/����.�X�����s���=�tm(��6��o���k��y�U?�&�A�D�|G�ӖK��\ޓ�� �4�]J�?���К.�M�.6���w� w�,~m~���~Vտ
�-�@�Q&�]E� M+7,]���T��|�A�Tv�P:3(5*��.Wݸ����o��A��V8���iiqc�FV��� o�0������ghk����C��6�"���i^(��0�ǋ ���Uٜ���4^>v�ƼP��";�+טc��@4��w�6�Rh;l<l�z��P
6U�W��O�ZՂr�+�;71��	�s����g*Y,�K�3O��:�BTm��}+H@���{�(�j�g��	�@��'3n��3���x
��v��Ǚ�F�-���4y�K{I�sv;X�`����U;�O]�ۍ�a;����N^<Xb�n0<djA89!c{���~Ih�9 �jNg��ځ�y;W����C��l�T�L��s�)�l��@��FY/�8�đ>��vM3�����N�w���Ŧ�2��O.�[�8]�'S#�dl��c6Ф��<��A0HJx<L�6��b����.������v�5�Ye7�
�a���Y�i/�,��h�j�2��0�Z��
��]���%C�41���`�&C�z�ӀV��\]}�=
j�׼*J���.���J�lj��׫��~-v�W�Sڟ,A�e��hI¼�����/���� �a��0>�^OPMR�1�m��?�S�U���̹N]|�Z��;sD/"�Wڲm�Y���6�P���2>n$)6��[]�*Ӏw�Bk&m<v�G����)��������]^���f;|���ޏ�x _��uMqä�z�5Z�80��Wp(6?�~�S1�aT��B��7��j/[OEk�M��8�
&��9ݫ�#�,Ȍ^�qq�%;�	��6t���!��(M����0n���t"7�Wc��'����"�`�W�T	@�uW�1����dj�/F[Z}��Ki�O2q���������f�5�.�+���k�K�I��vOM���9Z�B3���y�Y��ja�s��ŽXfS�����R�[$LKoc"բ��Ѹ�%��+�&V5��/�b
F��da���鍲�I�e���ʉ�1��V�߫�e�Ш�t�Z�� � �~��������#��J_��j}�[t�����ϥB�A��,%!�s	z�,����X�v�7r��s�`1����OR���4�p���uvGG�T��8� '��n-���<��5~됯�[BɉH�Gy,�R߶��I��T� ���|5���M�덽�+$b����*���)��ށR�3O	�U�.���Ѭٌ|�E�O�� �Տ��л��#���v �
.{���B;4�]�Z�<cL���5T�NQ@�>(�K�*]�!n�+k����3��L'��|��
�VT��h����"�Nl܀��`��ܪ��oܚ^er���B�4��m��÷Q�͸�h����ɏǑ1�o�	S2���&Oz��@�g���M�G�@_�iSǓ�b������Dۆ]�{n��hJ,�X&����Rˁ�h� I����h�l�5�%Y��H'yQ6�{1r�&��@ۿó��'�L�Oz���l�2����3�R��2v�W;Y�=P�	�Q�X�	-M_��fvQ��1��P�Cg2�Ѻ�ֶ�_�лo��!.p@����Q������>ݭ�O��2�\Ѥ\I� �;V^Ҭp�x��o(�4D���O|�~26���O�J��+��ю�b�R/؉�=ɠc������X�@(��Y�]��$�)1�	�(+D�.�?�]��=�4�O�zTy"A1%v>le	lo�����@�a[�a�����'v�==)\�S�Y�H����UxD�c0��{��	���1���p����E(�j�Q����F8����9	��O��[���ڂ��j5X�D��un�B�nF���� ��֏h�/v<sL�<4��C��Z޵-��3��X�1���[��ܼ��xϳ˩$�Aq��1)�:��̼D�G0%!�Ś�C����u&�������^^��0�p��^,�����ϻb;���Z)�	ʧl�PyBt�8��t�<TG�v}�c�IP��ڲ�+�|3�L�2w���zhaX��)���'�@���x��6�q9,���,IZ��܁	L�ҎW�.�xO1� �4"sE�;�1+�̎���79�_�@����_P����B͚��ce�\2e�SHr��*1�;��.-�m���7(o�����[��
�I]N&���,��F�p �#�`U9���0����sқ�;ڴ����t`Ex�Z2*^T"��]���,)��]-���#�;�]�f�=�o��`"Od8���|�Q�a�PJ����
A[0�t@�{)�J?�h�2�>~֋�}l۸Af�F�ʎ+@y�jI�j�E
W-�_�D�~L�ࣜtY#ќ�j�2�Z��gif��/~�>�ƞ�WN�r�('ƈb^�a�*bx#�#��ܹY�㳢�צ���1<y>e�,�'jR���Ͽ��cnV�u=N#�A�-�������ua��0#p��o^�C *�ZSkC�o�񹌌 ��۠�c2�����>&l�^�ƥ��2�zI��|=7�c(x�1X��^1�U������r�r��ܗQI�`ԩ6@;���~��[�p_�����0�8�9��m�ֲ{:�9��p�p���c���[ ��8�O��OuvJi���~�rؿ����_������4#�iI���Tv��:X��˴
��A�_eH�ᒴ�s�ӊv-�5d�Lc�?��I����^{� 9r��k�n��L����N[�ʩ��1��R��a�K M�e�h�u_W�V�1~��*w��~���"���".�	lK�
�#^I�;���z\�Sh�����C�EL�b�I�xW�����݆�B59�,��ә(Ɛ�qEƐ3'�8t,oĴܥ��sx
�4;f�S�r�u�7�`+��_�*<�<�1.F��m�j:���JN~��aU�6�,�	��c�7h1��Oj6��J�آ#쟋��*����U�3�6#: s��n�F��$z�yaX���"����I�B��3`����g���Y�<�KpM�x�2/3)�6o:�
�O�g%�{��i>ʍ5M���-e-���0@��2��6p����0[#�1�]��&���A~����7�q�M�����7��;#��,4)����чq$�=���I�%sxEC�0�fͅBO�B���O*Z�%0�	����6!�gVR�E�`Y��'�nhf�;Y���T
�W-]�'Qjl�2�oM<�e�a+6������J1�βt��D��Y��/�����t�صo쓝�G���7]���o\2^+(���i@��q��=nUO�y(�9�4.�X��y[_�\�r�jf��h��l�Ǹ�������v��ﶆ�E��m�H����
#P�=P��d�������D"�G��4[��DX�ax�j���W����I)��7 V�B��:�z1�*C��b�{[�+V��'�f�hfҗ�x(��}�`A��(�,BEUtkF'^?P�L���"Ns��v��Yk�x�⶚�����-� �S"�֘�4�� �����I! }����d��|N����.��������ٞV���ͤ���u�{{��jW� ȉ���|>m�aу��S��:�=:����ys�Ga�e�+�H7�!*h�"a�x����\��{����y&N���:K��R�%sٳ�l3��#H�� �'Į�X�r`-�z�ڮ�a�4��N|��rt���*Ѥ9*p��C�0���Ī��t.�!0>�E��[��5�:�oD���h��f(i����ĥ���).�5���{P�E|�bN~k�z��@�w����J�l
�=���'|�8Ӵ=_�t�e3J�!y�C�RUX_F����xv0������p�'V�c�7j9:�φg�YMK��pXǐ+�Z�/oPm`D� �(�������*g;�AʙDps�N�1_���'���}k�Ʈ�a�3���T����Jz�	'9�U7�v�����#m^Q�X�M\���a�g&7�R�+TY�P��vOu�;�%]�!� j��
@ſ��E�"W�!�K��4��(G瓂�fa��i��q�� ?*&�̫��>q6C��d�c�D�R�n,����V��T���O�A��=��ٹ��}b1e�w*}��.�OȹGo�94T$թ��w� {�՝��!��@�ƂgQ�Fʥ�ݣ���I�⡴�]�� ��?k�jA>�4%�슍wX8r���\�֕��Y�RI��)�� #M�ȼ�8p}��_Z�B��d$@Kj��C� dU��4� �q����;�.E���N�&URWD>��q�y�{��� Zp[�p��9KӘ����6%b�V�.=�a�hĠ�&��"�Sܭ�P�ݢˑ�E 1R���C�� ؖO��]v���1�AC�����;���e͍HC!��F��<;E��w D1���p*��z��-1A���X�:�<$���Q�)�#��D�7�Bl�pCa���'�}�s����!�ol��r�`�Dݰ5��J��,ME�7�����;g�(�VH���bU� d����$�D���.�������f�Q��xӨ���$�0��L"�2��W�v�,8i:��D�����a��c­���	9�0WȔAN�������S��9V,�/S�9�qx:= ���i"W�R��ߋ�m\αk=���.3��Nf�6���P�|�����!:;�.�����3��z� :��V;�l�O6��T"]�d����HV�KwO�?L���؃KY=��+��j��=���]�� 9�	��w�*�\;R���W�Wv�d�0{���f�YW��}&7>p���(u�g#�)B�p��sԀ:EиOl�<RL��ץ �������JP�P�� ��=�Hm�w�0�ľ���	��I����<3���ڣprk¸�a�d�b�=d��f�ט�%.(��2��Pu�c�`,���NI�3��D[�L�m״:a��DH�훕�p ɥ�D��KVL�V��~��0�=�w��z]�qC��n�Bx�߆H�?����V1>Sʞ�i�j\2C`󜏷|-3����[�SFס�pqt)8��}�'1-�^��Pة��%�H��|%f���|Oϟ���5F�� ͟�G~ͧ�=�p�M2x��[~������C�R�ŏ�5���|J`�m��#�8c��.��뭢Rʮ���@���2�q�ʖ��������}���G@%�/ro����`G�m���
+�o`�Z!;��DH��{y(�a�������}�.���.�� F<��rd{�>��R}Q�iI&����&����6oX@=o���e��zk�ajn�C�(��z��	�`iz���B�DxN����o.�7�#���L���r!��2��N�K�G�қc�n��Ӻ)>ꆊ0œ�ѭbY⪺	>����>\àI��|���b��p�p�� pn^k�Qӳ����_�u}�&x�ǲxMUFШ�;��G��?��'�gY�6��`�V�!~Ȟ�F��1�?� �c���l�*N�ͺ}�\�'�e��d�����{ +v��U@����u�6/��gd�RmCY�uMV{��Q��l�wX1�+M'��E.���.�r&:b���w:S��0G�
��=�a[��).�ű?7�5�L%��޲��?0�ĕO4	��Ki+���2)�\���[�?�ɺ����Z��Gi��բ��/�aR����<�0Ȗ�5��eg SdV�(2
k�%�^�JmP��/�� 3�B]m���?=���C�N�>{�K�<g�=)?�&��G�ޯ���l���̀�ʗܴ�͚�=3<@����r����Xv �8��|�^���2bgm
c�p�y� �&9Q+�y�5R��������:<[����l3"�u!�E�%-����(�{�"�Q��ֺ�{���c#�he�,^��e�]Q��wBn�>��º��{�=�i?M�`KE�	~6���MK���_1�d���Ps�ƞ[:�KC���t�֊���M�}��x��Ag4��������[��1�_k_y������o|=���d�'OYB��D1HB��C�u��(�������<}s1{��n��ԧ��~%O��T�KfL������V}1�v�����
#���H��s��� �☐�jB`����&!jή$���"�j	���=d�&��9��!=Λ�%"u�De�aOl�n�;�jm#�~�L�i����)Q�\故���B?1�T�p~���@ȇ栗��H:�0e~G��	'Ѩ��U�5��\������ț{�ي�6�Qf�k�U&T?[�4�k�(!6�~yвս�ܘ"�����c�����U�Ne�ڻ������e��z���1�z�qc.;7a�U*+)�,��h���48`3\���o�wh��Ļ-��������
F�W��btMI,��`�?}�<T���6��S�i���������+���tTԽ��'�o�\��4����:Pp�g�#�l�Z�q� ���ƀ�h'�Fb��jH�O��r�PqUT�1*�O,����:���kU�((V�.��[�q�G��Ǿ� �\�mm����ݝ_� U�ܞ�9T0�gX�,ę|�\�?U�tiP��U�H�bh����i�hB���@�'�N�yF�@��o���E���b˅O��1(.$�D�#���6�=Tv*�e�P�]+!��yH���o������k*����a?��0�4�\�L:0O��h�E�d������8?=m�850�yȮ���-�i'��/��������)겼.��~b&�KW��@���k��3d꥜�Q�`*Rԑ)>��R�"�A,�q��q����ܓ��e9SPd�S�,2Y����B����c'�h�֡��_t��@�p�S����9=i|b�\�����ի��_dLK��v�'�S7�����!��G�rx8��'A|�)?]^�����Z1.��ezy�|] O).<.��r ��:'��,�µ҉5��W��-=W��K� [%6ȰfK���|G�����P(\�8��{�O�lp�B�&�ז�5<1'z�l<���W�Lc����"_Y	�B:�i����p���Ĉ_�Y�S�ע���ROд���ͦ{��p៷6$
L�)I��9x%���c����4�P(��،��|tT�xԇ4{	.'�K����=K����b��pWƴo"P��ؚ�F���;�g�k�Ŭ��.�n�N5V�&�v0~�͸Q���BD ��W�J?���^�����>^��;�I���(�]��8	(��y�etw/Z-IFY�ui�����A�u�U�T���zoD��N_'W"�e;��tG����������	}yζ��uy�v^�ZD��e�\��+�'T�*�<;�'����z�\�Mpc��4:����p�8QUj���9*���ٚ�S���_�����Wj��s��aZ���Rk���!61�����{�V"����"D���T�yt]��֏���'�X&�p��29�fT�����ҡi͆��es/-g�ۢE��ȅ�n�;!�U'�	�Sv�z]�&��h"Cg����%�ʎ�?e��CQ-K��wPM�f3��e��}��=*x��2�R��9k���]$�^I�I[��a�.�%�^t)u�"�#L�K ��ę4qL�3�#��*�b�H�K���$��8�z@�� >�RI�]׷6��`<���%��o�xH����7�C��f ֋r-�5�/�n�M8@λ��޷��f�p���*E|�4�4����-t���ꮗ����g_5��gO��k���c��#��?ѣ^��!�.r{a�&���a>���3Ew�)z��*;A���c���QD��J��:2m����Q�� �(�U��b��;@���Ő޽���<����ؿ��m��W��SiP�?�5QXl�=�1^Ζt*�r&�L�Eƣ�����6&��r���MԝC�H]+����&;D8��<��m�`�����?L�6�r���%��-�mp�e���&2�b�����(���o�����6��\P�mg�L�Ɨ)$J���4�ʳ��-㎄n$r�8Sgj�|NѤ�ς����{={ge�[Qb�v3	�-�����.�ң�@B_�8T�	b�Ry�g?�&��:õ@�n�>�=zR$-������R�`�����#��}���8�4$ev	|-K��f՚i/�ڢz��L�[b���62l�a�hW�� �N���Z3����\l�aJ�mHn�ǉ�q�|�1vrM�O%)���c/q������\�_��f����=��k$�Cզ �[9��-���}��g���=��;�����E��#���D��b�,;����aY؟�Y\7���.Iq�Tz�G���D�L��j������ŧ:�-_٥ڂRɖ�pao�U�WS蟤��N�0��md(�w����HA�4eɷ�zL�σ)�͂���Z�-����%�>���4@-��uo1x8S���t�;��BaG����592�D�|�,Xv��g���':41���s�~ǵ�U6���;�
f�z�����8�v�%����\�~T`L8�6�l��>�Sԯ�ge�Y#�6��E� ���`۱M8[��K��3Pn{�����%Yw��5D�U�����o���C�)W<L������n�%'�;����6O�6��O�&1��B6d�[S+g�}�<<��$ŀ�f�'AX���&}����_ԅ�~�~tV�X�ǝ$A	*���p�A������J���B�v����~
�Qh���+�Ǔh��;En�㡜�waF �s�H�u��I;����U��9�R}���M5�ߕ	�H`P�y<6y>�<xk,d}	G}�}\����X+`���U����;�]����d����Q�M��m�x�D|��X�����{�<�8F�{�h\���F!6]U�7�����ҭOa�h���v�]�}�^gn5��	���R�!�E���+�E�����B>:Y��E�p�:%���`��N;����T�<ʒ��m)���	�/k=�mbQ+��a(G]��h{=+��׆^��:*֎�M��i��?�����!V��,8y��}�ޯ�?��a���_[��	���O����;M�;	��|��)�o����١F2�����NRⳊ/Aa�>#�ʞe�:@2�v�����
K6�"Y���,].�1]wo��Q����%Lږ�KmD�d���|N�����֢ts�]&3-R�a�-�("���o�M�:���mN�fĊ���Ṳ�8.���t�r��J;��f�W��~�7�8H�.�&��6��yZ*�P�D.� �����L�m_� ���;L���	t 1���1	){�^�c�e���qI7���q�3�8��QZ�X�>�K�	�X��N��i�l)6�%�1�y�������	�m; #�F0������PՒ��~��o�N�z�1!�^�en��~��Ot@�����۳��q�ILe)��@eʫ�xjCԘ�t
���Ȟrq������.mJ���C5l�KSN8�}�f8Y��p��N��yQ#���b)%��!-�
owJ�#^2|�N����1��z��v���\s���,� �p��?#���� ��0�k�)^f @WA}h^!pVR��FK.�%i���Tl���i��n�+��(��@=ө�E��Os!::S�J�j��vܜ��݇�T@o��o(�$E��~@�Wgk�� ����_�h���#bo��9-�Q�M�ݒ��%��q�+�Evp˰&$�B���sd���	�Mߎ���Gf䶃���&���OY<��$��u�K�|������؋%wڊ��'�[x��]4ܭu�Cm�A��Wk����d;�eM�,F+ �H�%�9|�w(?�Ǧd��{����;�؀�y�d��ǵ��%J�� ���H����ROM�Y�T U}�ܷݷB{#��0m-p�T~���"�B=z�dڱhb�% 
���!M��3<�� �F?�8����p�̿⇒�EG�){Zs�6��㑨p����e���<\��HX��(�EVv�SD� BQ"��N{"}r�쐻�fwï��X���^�*"��7(�I�x��2G���w��>8�*I�N����ʄ�oH5��UR��-? ��P3�e�
`��X�oh��$�b��#y���y��t"���xh~j�EW�0^c ���"V�&�X�rp�M`� d��SRZh,�;D���/�ᑏՕ�s2aw~�m�p]U�Q�(�S����dm��u��l>a��^5拏WzԦj\��P�RaE�����)Z���YW�)n
��>Me_�����M�uAd�
W;̓��;84|���z��.�v|]����		���Ʀ3z��_�D��f->]!v���,�*}<��۽�3N�#m#rp��w�5�/���q�Bct����l �7����}�b,b,ݐw|��2��7	�Co��u���cn�bI�oZ��$V%���t�S��t�JI=�`��zI�`e��U�3籉�+��ZY���!�N@Y�8�e�׎�BF�@��с�NU<^��ݞ;��N(�t�l9�~�\[�|� �u1��q�q��,�[�2��?M��'�4�y{���L!T��r&6�$�$u�*�3���u���)��E�z �k���%�6��gK�t�	�B"��v��������K͊��?��(��BHǇR�D1�Fqc!c�M���'�^����؈�S� ��mɰ�a��)[p`D)�#%n o	>��;�$����E���ؾ2֛7������Ni0i�s���~�sw1�Y��хPDmrH�rĘ�t�h稧�(.���b?���`�z�_���I�X��G�5tfX7w��ˆ����F�zY���凖�P���S�3�O��M]͆�t#�k�Z;JM[ �U�B�仔+�B	���CD����J��S�6��7�8�$�<�����/6�Q�f��G��b�r+�'T�ស�d�ƐUq�=8����Ȗ���`� ��!h��|1����jN,)g�3��gT`� ����N���x����n�07a
Х*����q,��BrqX��~�������GI�[�������K�����M�j�v�f��:�MCG+����ο.�5C�/l!��cvv�?~W��b��i���y����Ơ_�E����w�:�eH�ƶBQ���~2e|ܦIb�����T�sҼuȢ_yk9���|n T"͑"�M�@���,�_;�p��#�=yYS6����j�\U��r��1K�LU&�;��7J4X{9�b�M�Mhx����%��Y��M�Ks�yq۴�(����Jd&��i�H��%��ࣄJ�$yQ�}yGW4j��.k�!�1!6�^N�o���CLӲ�ɣC��	��2�����e����2���!BL�3��ݔ��r#�}��@Ic'_�yS�|����y]�f��	n�KʁSL ��=<�Wn��H:�� ��ؚD<Zݨu0
�.��\$C40�s��.��d�5��tY8F��^��Ul��&��Ud��rCq-A�g4/yH@q�o*J`�%W��T&A�F�Е�����B�ۤSE����yt�!���d���3
6y�:l�^h��w��*)@Zk��K;J'��K=!y�ym����)�+�3��7I��q�KBK��� 5QZ;ᒂًV�>ؤ�s!�rg�ՠի�,��B���nb�[��+����)'�\��u5j,3>�.l������iO��t�;��X�K���P"8���=C,)h�Li�����&@p���4�9����u5��b7��K���P~48A�/��v��$<�P��[�_��� �R�P��ϩ4���L�(,=�=-ifN���V��Ŝ�p�����*�ȗ��URI�^�.��&3p��][�s�?Eɱ]h�I��l�y���I��?�[��<��6�fѲ����{;/.爆;��l9�J����Z��԰�lz�I�ŝp�E����䦤�,�8l�\!��K�/��AC�%h�QҶ��$���K��x�����;q��֊�%��A$���$��y,6�� �EG��D��tc|��ؾ$���:�!�㸬5��<�j��	6dE����6��%2����v�y�)ts{ȟ�Y��=-	�d���W/�i3�����՝�e��מ̪G"�*
�]U�i]+bOsbb���pW��+�/���Ia��>�%h�����<3BIz~��D�%'���2#3�Q����6��L����ٮ}��N�
!<�|/ϡ�@��:K���ٳX;�2���Xp��W�Ϻ�+=�ۄ7C9�
�%>P2����D@������(����j��@�41l	��FE}����}k�&��Xt'�\
�R����(\O �!�B9�m�Y[,1#�z����mպ�y�ck���p|�f�S<�����u���1:����ņ>"[�H�n���0�z���]x?yY�_3X��'m�
���}3�䶶��,舃�W��٫��oiw�Q�IG��h2@s�Sq�ܚ��S��2�R9G���*]{g�f�$��T�*t�phrW��Ss�\�'W������F�T��O!�B?�!D¯"�1�EؿP��.M�/x��H�M��9�<��k�|�"��Z�-�:gRl�I�ʩG�Xȉ{g�̤X������x	��6�i����-�ٚC��o�^���>��^���9����R�~�D�����D2�A>5�_:w�7- �·|�����p^�^��<�꣭V��E;��`&���N�,���S����O�%}�_V�H���"�|�B��!�'!ɕ�f0�z�P�­G�#�A�#�><U1�H���������.2�e �;vn�9cL�֋ c�7�w)�;�Z���6�(Y &;�,�
w�g`0�ϔ��fHbN�VB2u4D#ʲ�c�K=�}���\i�x�^����'f��%�f����^��p���y��ۼ�IK�WB��E�����/��˻�p�Js��unт_����pv�Y���!�Y��P��9���S#�h9pE6�N�ͻd�����;-�� 1`��LT�{�9R'lQ'����ӆ^o�0,���Q�fY:�.��v�:����t��>��P��꾲�R{G /�b�ha'<�	�7�F�7��E]M�\i};$  �٬:%;���k��o��}�w��Cd��ҁU�=���l)�9��V"�[���S��vC4 \�t��?��h��e�^��g�G�ߣ�{'�Iӈ�Y�+ĺ�>�G��`{+��{u�Z�C���ѽ�[p�Ra�G���e���{�X��A	]�No0����`��`�潔N��#�����B���u���vJy�[r�&���¼h�õ���[O��� ��IKZ��T���� ��n<L�2"
Wڴ/Rx�,�ܞ���g���x�DW2��48��9��Ƒ�ot?�%�.G�̀ňC����!��꼶�w{Q]�P��/#W�]�����Ԇj���s��8�ۭa���J��F��H���%���[�\E|�ީ�){C`��M�(F�YR��B^&�":քe�L\����NA?���T�0c��~I|��!�?�i��>��x�PԬ>r���l����yt��D��Cy�	���] A2��$Kf�p�ɽ������ݮ߾_ru���$�D�?V^Gǌ��z�����c�4*(�-~�a�ڛ<k��)�{�jx$L�+��?�]VW�br4�}�Oq|W�Mw�`��������dH��VLb��֒Ŝ��s�(H�e�����0��0֤��쾑���Xq*��r� |z��T,w,]&W�V{k-�k��
�!}�s@�
8ƴ��P��FE,���Qr�ͪ�Ũ�ƪ�Юk�mɬ��k�����M���Fs�N��;"(X#��L[-\PvȈ���`�E������r-t8��ɻ���_��޴����i�l�͔'�LW@/���a��Y�5��(�v���ѩ��4Cv�^��:.��N���#�a0���E���g���PS $�7�&v��UF�� D���Lj:+vM�{�Nzg���5b(K��Ŕ��mD�7fO����d�(;>�Pf=qz���J%'^�tH���ޙ�Y<�)5���F��8�.����N�vN|g֨"�ϡ;r7��If��Ǎn֌r\u�і�(���:�ؼ�ݗ*=��E��7�	�g�^�	��Oq9���I�*{s�R�v�qۿ�n���e���Na�ո��H=F����
i��2s��䛢�ITEϽ������QȦ�L
1���F3���*�N��D�6:�� ��f�i������DGY9]HsʖS�D�\�*��p�)�����Y�sVV{���K�ٰN2��\B�!L�/tB�]��c�f��Ӎc�!��^9�C�\Z����w�%�B�� �RF.L���g&�08��O�i�93������W<0�x�/��R�s�O8-E���mne��ap�:�9p��=\m2p�=���ZL!��b�@	>���j��g��(��ڃ�K��e뙀�f4�`}R~%x��KQ]�-M����?)�f>�1'�lI�5|�������>-���)3�
����(+���n��?H�|���:sCs	sc�*<�T=X::��O�k �)�[���Q8%�x0&
[�"���.��5O�/X�#�^���	���~$?�еEg�JG�d3L'����U��ҍpg<�w��<��5[W�2Q�V��YRnG���8\��9�M=4 9���� 	]+�FK��-�a#� Zܜo���r�J�.�O?n}�Y���K�3PU�q;Xlxc]�r2�̢�e��D/Y}6m�Bu������ysȲI��w҉mhq��� hn}�ZE���E���Y)����m(�W��Vhg�{����3���6��JA�)��|��E��9�\.�;TԒ�Sb8��\���'�BtE� �)�_2�|a^�ضGf!�v;3�{�-�@C͡qra:)W����+���[n�r���y�餉��M�Lg[]Z��u�l����FD������(���C���¢v��Z`�Jֶ�C�P�]J#I��W!Õ��1�;��	�pa*/�G/�`�)�8CQ[ND��Kǋde<o�R�>#��M�Drج�|��.�?;Ͷի��t����ou�F�� ��UUJt�ةFZ�����o��=����kO�r0��p�S~Gؾ�"M("�.^��Ʈ����O�F��=��!aՂ�N��'9Rg��F���!+��Yod��i��r�E��kyN�S�b��azU+5���n�h�k#Rz����qK�	W��$�W��9����g-�O�q���6A�t��U�b�/�v3`Z�c@}�̷�I}�K�l���`�^V]��=X���`�]Y��v;�/�ې���(=c�Uhs���_�)������&����v{D�X�YL��n'�+О����\����)	Ձ����b�|�V6W����3�,#��@�`���x>��T�k&;dˡ��ã���}u�
-�udq��̠+(��"�yv��sm(�x�5�yD���~헫@�>����yKW�pw0�娿|PR'CY�0a�#�S�p#mD��&����rw��J_3���g�)*��K>:�!�� j�c	@�Hʖ�7%)���g�oh�W&�0��_����/%S�Q����c'�+V��+:���Mkq�r��6�1=��������뤓�*��~6}/:��ɑ����Z�� .�����J|h��*pϞ��E(�A�g%�[s�6>��*��i!�`#��k&uߞ��]B�=�O���4.P��u�1�׍v���yy:�w�K�8���x1�.�k`�M b]y3��Ű��M�K� IP��#�L�}��A���Pz��_�_;�L��Q4�{�Q���V-S��b���߲Ξr��~{�
�0�Kr��l���/%��
Bpd����a�ή6�IW�
WfN6�y�p5ˈV�hH\��!g�8��p��;����S�c��b����W)�l�Q�GV�J�R=� ӋS�xQl��8"$��g�B�[����!��&��o���*x:Pmr�������sv&^-�U�%�U�T�r*��'9 �-7 Bv������(ؼ1��S�w+ܫ��p�	���w�����eF�@t4Q�k6��yza�t��]��^/����|`ҁ�h�^�N���
�S7���?���,w��f��H�p)wV5<��elڰx,��,�JxAB$h�����붙[7�ըV+��0D��I���I�v�R��<�^fb��H<0uO�a�J�Ш��4<���_n�1)�F\;wQO�S�ł�P��|�~�>��!x{o�Nd1\�l���!^�k���6�%t����G�4ԢH�\��]��'H����j���hS�&apk9:���j�z��!��@� �g��Y���x4��Qy��K��A�����>n�;��%_D`(�1������1�vה�K�Ii��y�`�"�&8�&h�~$ܧ1,d�9>�`�piI��"^s��9�2�w�C���IE��uϳ90ڣ�f�|�i��O�(���鿴!��4h�f��V�_�� �Ϥ�٠��5�x�T'e�7_���KB���2����>���%��z;���ݰ�J,�l����B&�F.�r��g�Oݖr��с^��ɼ�(V��ё�X�kR��`?Z!�ҜHʇ�������1lQC����Hh�P���j_��dǬ�{dbK��]_�I�_b�Ƙ>}��/<-o:l���1"��B[J0���&���t�;P��;3�3M!K���}%�n`")3:R�e���݊R�僃�;�L��_���!yᗶ>�t�I��7�:Y�$i𻪕�f�-��!ʧ�V�yW�����1���C��C���}z�˥STZ�M�Vtc���L�N*;�����\ �:�ݽrw����P��!F@�r��ʓ�y�m�h� t;�`��6"y��s��`��:;w\u�i=�]�����2�ە���:M��QX����o���Ůïv?��`�n��͘/S���_c�}� \؊��{�A��(���&z��:9�/~�![fɺ���:[xE���Rf�q�6՚g�Ȯ� ɩ�iN��ܜ�z�F�P@s�<���)�_�Y�O����Y��iOMH!�|��#`�Q���������xU�^�}tk�xj�����3����p,�`��_�~/t�FZm���p	���7H���Do#H�   U��_r̎ȣ�"�ʼ�;h52z��sI?�YY��V�-h�e��%���1�ѥ�����F��&�P���:]��Qr���&���nF�F�_*�c����R�z��#Z�#�&Aά�ZJ?2�ʦ�s/x�eb����ۅ�qoY~bU���9O������[���x��\��L��&�T����e��v�㗇��5���*�!���RDK��2|��jƬ��VF<�|��8A���.���:�cD��w�2�j�!:��C��^_|���7�" ��-e�+&C����������6o�ۢE�o��H�Ҭ��,v,w�[�;�_1�gu�ca ��M)s������t�n�!�'/� �G��MRY祐*,�i��e�:Y���b�Ϝ�h(�u��<E7���9�`Kk���8\L
���o$#8���B�J��8�� ��x�Lߝ�����\E.V�{X�;[�tO�ߍ$Ze����}m0����<- ����/ 6d���!���c����'(H���ƣ���݄f�o�����x�w��5���e���]{b�o'�q�on(����JjC[/��#<��M�V�V����X�g=���H��(��ˤ������*��mR�� ���������)�:�bx���V�p9V��r������Z��L�s "_*��W�y�K��&�1=z��2��h�G�@�E/���|�Q���p&��rPh2W���5�-�iK��v�Y�vus��]���3/�kg@׃�����V��e��\�[�l�wR��#UϥFb,a���K���Z������ �\�'���}��enn�iM�*$�=J����U>��Q�8s��t�v�?&S���G8�?1�ף,Y����W�3@%f7��N�x(q���rJ���(g�䀲a�Ѓu�J��G� #���UF��:۽ZY����o�HMd@*�:[9�M�J��n4�M�:��$6���u�9�(x��ݻ��Cl8m=+�@4�*��!���+�>��n�=�����b!�"�~BS�\O�K/�=�.z�0�{Z���_-w�(�T:��F:��QC��MR+O�߆��7!�����ٰ�H�TA��$ht�=�3�O� hQ�7q%��JG��IdU2I�����8*>���s�;U��N�)��?p�e��0f!8<L�,Y)��6��Ѣh����e&��c��%���Y�o��8��:����j�6�P�k��Ƞ�4�	X*��������g�%f2�*�BF��D;	��Sa�)�c�L��`{H�c�.�R�� 佛�7���cj�yd���{�v#���;
���'!H��4$������硱�u愱Nsܵ��M� Mr�(�j,�r�P�m�9���o�r$~,�3~����,� �^K���Iy�5.��<x���6H�G��m���u�l��p.��%x�[�̰��1a!8R������h��Y��z��)�q^$�kgu����p>T

�}&����JdwL���{!��7�82���8�����BH  x�Ԫ�i�Y��J�:[B�k�mC�X���M�m$�|�_��φ��e�b�lޞg7�՛�T��
�ґ&_�훤o"��N/�j^��BW�6u�f�*��o�6_�`i�&���*Z��8V9u�ր���pQf��)" ��3���lB�b�C,�)輘�,K��4�X`���WR��0<x|��&�����}��"��LU]�̞[�}�l�OlV�Q�DXb)��L\N��q���3][]׿�@�m��^N�#W#糠��v�g���4v�?P#ßn�4f��-�G�?/���m��Dď^k��PeD���U�RT���������ġ�Z�g
V�=�ȥ�6��f'v�x���tx��W}P4,b^O��qDΨ�F�7��L�� ��&GY�1X�nM>aA�L׳�U�����/�����u���Pu,���,G��ȝf  ���B�@i��g��#�@q�WIA����e\&Ʊi�{�+�R����J��03]V����%�SD8>23����oȫ;ͱ���[�sr�~�z���&���`��*�= �� E��!M�嗧��0Z���"�b�}c�U�)����@�G�g[`�O1��]�Lu ��ar.xR|��&�ԡ`����D��-Y~�,����~�A�Z�rP�{&@W�~��u��%O��,�f�q�[s�N��oJ�T�=-�?����լg,�n(�޺����P7@��`�gM�E����o�����.�O��f 	\���DdD�Y<�\��3�!�/�_|=�0����!\#7���"-\�F���l&%ֲb�?��n&�~1>rf��N���O��O9������W�ІX^X����o35���٫=�;�}`;����` o�hZ�	Z�$ Ы�>�l�u%�k��K�֏��^+��Ŋ�o��3�fdV�|��	֝��rl���Y�Ę�-��^[���v����[�2�W/������'�)�'T��E~Ý$��CE�h�=Ϫ䶜v��Ϝ���o�c&�I5Q�|�^�bo�м�;���mޡ�ͺC�pͿ|��
I�d��i�Ә�d~*�`w�&����X����H�p�4�8��b�x�-r���%ǂ@t���n���Ԯ�A���=Y?!����K-<��n�rm�Ti���%1�c��%jy֋�3N����sYb9alda�\�!�dn�x0"a��^.|ܥ8&�W���Me���3I;�)�zu���j_88D������[�b�"n����r	�0XЫ3�ù+dK��w!��|�V��Pa���P���a;���ml#��K��xNq;�8�UN��!�{a
RQ�\�H�e9��ݓ�7�`�h�n�aO\�u�
�;J&>V�)��v!�&H��`�#�˼+FX�b��(H���k3F��4r@ Y?�%���#+���
x��놁{�!{�|�%M�vԞϨ/|�m��.(iu�n^^�|&��Qk8���"+obW��x�T˙���t���{�~C�Pl��S��8$�kfk`#���� �l�fV��wgN�N��:C��.[|Q{)E���g�D�ɾ���X�a��4ܮ�5�ڞ�����L�H��嗿*�Q\��>>�����zE��@�oJ1�JH���9\z�CIG��˪+���	h�Ť�r�׺3s����4j���߶�4�2�7�����N&�L�;k��C�؍��z�W�JE?q�STs�,i�VXoM��=`@g��X�=���� M��=���;����8��(�12�}��$��lm�e<%�U
Q���rά. ou����B���[�I.���K؋������lGאR�'���l�Fs���6. ��f���0�ޠ�,� ��w��k���i��,��9�W�||7�����Ѩ�T�7?Ĝ��6��DKo��w�F}�R~c#�)|��Z��>f���.���{^?�� {,�-T{d7)F)����읐�D_U-'/D2�xf\�q�&��ӷ�J�W�n4��-�O{���t�����F��{&/`�_D`��B�'TH��