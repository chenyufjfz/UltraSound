library verilog;
use verilog.vl_types.all;
entity test_ultrasound is
end test_ultrasound;
