��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�z�b�&��R�'�F92īQ�-��r���n�]�9}:���=YJ��N|� e��3�
F2��w�*�3���� 2���1h?�vˀ�m,0��ZR׻Q��Ѧ�l<뉈���[g�Ђ�JR�M�I������?ON�j+����=*ߵ6;w&��A:��^��=:�8)���/�xʼ}!�Fʄ������F�X�E�̈<�L���&'���R���-�ԫ�y�(�oV
��Ӑ�G�1g>Ъ����۾� v�(�|ٓj�F~UX�|TX�}�K��p�A:���	��n��������I�[��|kSI sT^!\]�����;�L�F��t�/u(���������#©g���oդb��x��)���ڼ!�p�P��˚��[
�)I�Y:5=����v-0������
��B�����%�����{�� �fi���m(W'
X��7p�kl=CݵU�n�ԝC�A4ɕ9�{ȋ�ʜ(��}Pv_ ������
� -�/��S�r��.��I�F��v��Ii�J2�G	�?(O�kՍl�t!���A�A���!����&�N���ώt
��9;��w��H��5���E^��R�����Դv�8� �`�W'#�K�׳g��$��tT�-��)��?{�p�
I4	o[X��͟ӿ���|N`L"֧ԛZ�H��N���h��u����KP��w�urX��=nM�
�70/���Ԟ�`�$Ҩ潥ʎ�ة�	C�"�V�-�1�.@G~�ؕQ0�d�-?肁��_K��7%�|K�*��8>�/�S}M�Kֹ�!?��=^�� ����ފ.i��d���<vh�3�V�z�,S�>	�@:� ��{%$���|�1d��q���>ΧŔ�;X+P�q��<��4C���~_
'38����<wL��3�����h��:��n�-*0b��
�B�曟Ќ��u�i�뤏�@�x03�3��Vۭ�SQ�ڇ	�dEG�S�J�N�j�|�M�F߀�����������ĹRW�}�S��L�ΐ�C����7&ׇ?V>}f��<�k	�S�R} �N0MEU]ĢI�}B�P�6����4����h��(@�;Š_�C����3P�8����Wl�y�3�H���E-'O�	��!���h7YK�Z$�Q�ܙeb;��Pu��'w��ꞧǛ�? ��e1�f[~8��h�M�wpT �,]$���N��=�5*�.5�ґm�?�N��X�|w)��L�4�:���� ���؊Ac��Ƌ�}=TC�g��jl�0}���֮G��%��#�]qY�m5��7qGE&Xx"��t��N�	����\��  �#��M�&�,)��*X�Hx��_ƃ>x�X��9��Kl�7l����۳��TN ��]`��K���L��R�8Fm�数��%���&��,ґ}{�8�L����.�t��AQ_'��m�� ���C�����JT�^D�29+AK�\�Ӝ�dgo{�Ϸp�+�v�Y�-S["D.�c�E����1b?����0"���Ff�xR-��_�3o�Ji�;h4#�nm��j>�?~�>2��޲��Yt$�7ȁ��ma�k����R<6�t-qn�+,�p{wK�s�T���}-YtLu���K�YM�ƿ��M����$�c_:���Ԋ�v����^�xF/��e��)aJ����&uz�xߵ��-�H��l�+J����R����E�ք�o��ӻ"�{�!���X~�1W�_B5ř$F��G&I"���b�pĉW�W99$1��n<�a]=�^���a|dR���4�r��&�JAأ�Q�ʣ_(�ܒ��9��L&_l���	�^Վ�_3�6&�ﴪ�L�|�vG�KG�0E���?��I�����+�2XЭg�0�7י{�.~ ���߁���L�V�4𿊓����%<�{��>f ٌ�e1�-��p
���Κ�����f z��#�X�VG���K�`��>A�j;B��˝��
�ɵ@�T��q\�:z����������� ���s��Ԫ�j��Y"��rS\�����ID���.-�	��C�"_��{�s+d��$��|UTv�Yu���2sj��ġZ��e��EC�D1y��
-�?ý�!=��b��lT9R�	7�@O;�|�&�;\V㖌p����D�Ƅ�oث��=�ܽ���?��5M�ռ>�ӡhh����O�,~�r���ǼcE�P@�%d_D�9�Tt��Z�}~��g����r����?ooN�T���D	A�RR��5�	��Y'�M$�6������zҨ1L�c㯀zãg�\E\�����g���4C����+�<�+��"�p�nJ�,���Q�=�J�	��]�e3��L�N��&�8���-o\}�q����}:�?a�|�ŏ��T��!��JOfp�W[di�5�Q闬ڎ��񑋈�hQ�z��������Л��(��DO��Wx`���*F������ox��g�ܡx�h硳묰X�b��[�5��"��GL�󻼐����/����S�1��� �+��8�Nz̶�=z��P^jqG�z)��Z�3d���� �C�罍�v����8��	��޲^z��ԫ�=��;2�����M�C�}6��p-�>��s=a|����&�X��V��no#�:i;���1zl�(���h��#2G9,*�1�Q��ϥ�MjTjb��׆�3�S�<���Z���g�qŀ'�ڌ]�>�|<�u�[u�i�F������V�E)َ�MrT�~[�ګ3o}ㆨ�p�薮����)P	_�� �9�T����RB���l"��&bhON��=��(�Ix������*5n(�vgv Sj�rZ�&6��Z�)���CjM�����pn�t�}˚����x �������'!�������T�wAbD�����5���J�GAB Aj�ĸ@�H�yl�s~�ĕt�0�@�}6����`mFg0���;��� ~hz��-"��6�O�/[� ��r3u=�����K� V�s~�틕9~����N]y�𛗏���	U�%u�[V����Aa��橃����.�I����r��l}&���̈�&�nx� �y�	n]5��K��� 2����X?�V�˄����3[]֑jvf�<�S:oW���5#	K�CS��`ֆ��>	��IMXm	x����ݹIWKՕH�4�[Ɓ��Juo��{8h`�Q�@�K�DFڬ��-%a��_!���A��*D��kN攻�oV&&O�.��{�m`=I�� �˄w����׫8���ӏ[�����׆�L