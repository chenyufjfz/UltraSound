��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+e�ҿĥ��L�.R�d��HH�~����1^^�]-��s�T;υ_�� g|�H�\��#}J�� ����BW��m��3����"��8y	��/ιN��fxΈu��oo��iD�Q�u|��:!�!B�N��֜�x�]Si�R���{pm��k��%��?�~v�F��.���~�m1x��<��ͽ�Q�ҁ�Cs,;d��p4\�7�O���y�UB���δ��7�AGG,�ˌ��0Zo����\��y7��iC	��O��B�֩���2��Vz _����b/�K����?�1��k#�8>�֯���:�P(�������<������ ����j,�-�z�#�I\9��Ġ�&����?�ύ����oq��?Z��P�2x�� >��]Q�X7�܏|�� ��p�)����	^		,U�����zO~�͝��5��*�E~�yNω���=��D��fJ�ao��5�3�w2��*�����0	�Ds��E�!�\���Z�'��%ɚK�/�@�ue9d�2�
6�g��"���4K��&�ܚDg�*,�
�''c,��a�6V�W����}�<��w���4���k��x�^�|����^�Y&}�܅�;��!���s�Q�YЁk�W�W�f'/�v��͐Z��
�h�~YVZ���[�E&�d�Ep�dv�Zv+��A5�HJ��{��K�3@��pZak��#K���Rx���S��߀�j�T��+Z�7чR�UH8�@`6 �#��˅�K������4l�0(�`k396~p�>�IIkM�q����s���>,c���9w�����Kc�A+[��oC��jٽuLk����9'~6^q����-R��C/��������%!��P(��:!QP����rw\�)@sEg
e5��8�5v�d �"8k���(����Hh0��(�-p4:�ٌ�K1~�~�W��Q��s.�[�h�����@9�5��
�풫����'�4ԭ�2 ���j�1����S��A��/��]�(
�ͯ��B �������X]l��~�-/q��������vg�b�N$m��p|s�z�uK���ȖϞsS�%sn0��Wjc���b���͐ZnF] ���;ڄ�ņA��d)݆1+��(t�����N��ER��D��{-f�m�j̒�+��e�?�1�̤�'Ę�;��JM�Ah<�l�$�	]�2��Ɇ�LE�����B��5HYs`,KG����\e�ExM�fh	ן���އ^�Id�Ь@�M[�-��`̪��`]ëJ�I9�ƌ�ﬧ��[|�TF�_�w\�&A�������;4j6+��!�N���t'۪�����T	F���b�3�s����Y4h��������}av=[�w�!��n�nd.�M���� �H� .@0�G0墷gY]g�����i;�g�1L���"B�
E�����9��N�z��==����K�Aii����=��NuH�?��+�Mi���bK&
Xm�TO�mY2��2�����"��W9�v��+@3���ޙ�|�ù7ia�B��<�O�r$2=�1�a����{duO}Oz_/
��X���0��W0I�SK�3�Wp �y�έ�}�N��=�T?܈g �t@�M''��T*�Ü���Jg�3���'�G]�h���V�����6��޼�b�U�4��+,���J�u��6ޑ$�����nh���P~l������X�-�Dm�P9��6���h�O�j��Y�SG��T�J��a����9��܍z��������ɔ�u����͸�.�ʍX^�"��P��c��-�umԩ�J4�Tb�}c�׉u�p-��:���m����������(���>��^�u���cڛ~4o���Y��������1�-�G�%IzZ���C{�ӹQ�~��K�(o�>Q�ŉ��9��+L��Ew:�^W��S��J�~I	�rx<u�Μ�n��Z�3,W$� C>V�G��ɼ��Lir\7��]?���W��L�Č���I������l5�|��]܃���qYeS�A�a�)�uI�Mo`�O�X	U"�
}@� Ͳ 1Y(�m�.ZDb�'���:�2�
]�(��9�T�՝�O�u5.}3��ڻ�9�����cR+:,�w��^�K���}W����}A0д�3�*@�{��wc��ige?�<Q��֍2���Y,����²�Y�������������Ѐ0�J���n�9�� �c�&�d:ٔE��Pc-��9�3,��!�9��g���!n�(�M��2��ōm�,�է�*��C�,��$���+խðԝ}��J%;���쒵��r�S��cm��6<4�Z�[����bZ�QP����-P��ٛ%[��:A���O$`^86#��ٛ�~pqݏhU��c���ߙt"�j�\���`�d�x��l+͒�i�.��bQ>�[7���k;�U"a��PEh�Y��2�s�:��f�ta#�!���4�I@/U��eL���~�~'���92=�q�K�&J\f�sƚ,@��F�8#��d
˽�.ἕ%ж�Sq�D�nHب1�YZP��$M�2�m�R��Κ%gH=<�J\;$�>� ڰ�u���0���5�i�ElZr1]U1�H�I�D��Η��9�����5�H-�L�2m�(z98̫|aG	�Yd1�(�$\hX�G���{�i�
��p���M+b������'Ea�̥�i�a�9��P�	t��bMY�>����>S�Z�G#��u��؃Ʋ㭐g�zXpq�?��C�����g/�Kl�!k��wP{�(�k)j3���I����J�tD WP�ߖ:�6 DI��N����\T��m�RC�'���{����L�<��5X�e�-���*Դ��2\��B�{x&MU��t`8�����T-w'W-�`�)��X$۪eƼ=�}*{(��<������B+ �,�	g�*H9:��x�ꖱ�x����G:���<���L�r�߻��zN �׹e�e��w0�s1^y�9���Mv0�_�mO9�rL����g�V�ڿ��M��4�� ��)hkHW��m	�+ ���)6u���������Y^���˺�<���'1
��Og�hz�9o�)���wjy���f���ۖ���ʕ�(�Gx[�Y�E^U\��BM|��ԯ�uu\���C?{������Hv�0g3�������=�*�ڕ��s�A���p����+���KX!��`�+(L��T��-���s��>,FE(�@�]͏щ��<C�5��뮕��Ȥ6κ|���a�KF[��rC�yvT��.j��D��j4S� w���؟L�%|Ls+4���[7��Ȉ��E��t��l�1��r���j\*�������3������b�G٠Wf��e��a6^�[���T�x����4>�@�f�[;���Q�&�պbn��G=���i(zYM��?����c;Qz����Q�T��?��u7:�g�!KN�$N�slU�yN��z�E���̅�_T����%yHeJ�T@�����c�|�Xh��ߥ��,���	d����_G�� �Q�y�(�Gr��qI3�yPV��Nf#a/;C�hEI������ϦH�Z52Ě�D�u��Nbz������݅�C�;����gB����\.@ԕ���� �]lip���M1���}�uH�ФJ���b1��>Ã�}�nXț汄6�M96�e���[����1&��Ԩ���u������tj�A/d&��_��DL�)6s��#���x������ߟ��Է�J�g��;MvN���A�����@K���Ӓ4�E�2L�S'D����,єL��X�+}?3�y�q	+E["Cr/v0}��2��dSY�Zef�)z٩�}�P���������̮�l�H�i���|����T�S�������oiֵ���ۂ��,Vr9�,%G�b���̙YVyN�R2g��z�A]�χ�I/�������ȸX��qLL�{(�)�E���h�]��GIY�_ gü��C	�Fl�fZ���"��ꫨ;���1޽��-�)����r�t S�f�?��38=�b��{�5ali�ZZ��$kg�d��2��'z�c�;x��S~0�j"u�����D��cA4[��!�V$i�@�j��v&M��iy��*s�y������=�,[�$���u�<�p;A>i��%$`�����C��ҭ
D���I]�L���]	�al���o�b�o�ٍ%B��`�L!�c/��ًo�)�)8;ٍ�QS�j���H�n���.�B=g�Ě�{?:a��s�K��r�6R����w�1�f����$�F�<e�C_�>���R�r� �(��a��d�A���w-T�ᤁq�� �v:��`���zu|d��e��4׾um�!/N�����v�F���gy����i��M�)%P��$���������� !N�X�G
�~���$�P�ޚy:�~��08q7[V��j��Q.��8���o ?�(>w+�촿@'��b����q6�
���g��,�4�U�5�ʇ=򭮱%��U��	��XX^�m�>F�w�3���j�Õ(�I���Z����Ƽ_0�:_A�a�j�܁�������u�6<+�u���*r�g�"	|'���3 ����E��8}SuN�N㤧�M�����C�[7<w�JdA[h�+�I}�2;�e��]�XpB������ �����c��:<2�$$�*O�;<��r�Ն��.���+�9�z^^S���FԾ��Af�}ur>)�J�	��܂���}`�����Ψ,�	r�eR;�D���a��o|��D՛BA{�#���}���	��D7�D ao$�ʲ2��k�Ȝ@'rc�Y�����-x�c�� ��f/���l��:č�@����C�g��9�y̾L��zH8�?
�jQ	��Y1��I�$�Iѫ}�����2<2ɨJ���ğ�θ��v�|�C���P�"Wf,D�2Ssbf̙ҟ�3�iC{NP�&�"����|I ��)(L�d>x[����{FO�&�=�`������y��LǦ�������r�='K�afN����	��'`0z�����O����|;r�!���o%H}d,����=;�R�H���
Zp�q0�6�VWjj�l�v�(����Qm؅~6K���)�'ۼ���j����B^&��̄+�X�葝���A�ñ�쩝)�,2����p7:�lq��]�irVc�����q����K�F#[�=�M+i�����o8��ɝ�ݫn˒v>ޥ�������Ő����]I^8�'�9�j�א�x&滶�1��㲹�sV'R���(�@&醁k(si\)�=�_��
fDko�,��LX���ɵ%I�7�!R�#�~7�9S�X�?,>�$�9���4f�H����c��}m%��h��XԠ��1��r�Z.�: q��e�0��	��z ��{���=- ��z���ィ��s[���U��~j��x/�<i>��B�߼�ݙ!bY���ͧ�����+
��=&d����"Hw�iZ�؆�I�u�;hٕ��|�1=H��ԉ�ۦnF� ��0l��3h����
�Z����:F�(�: ]Sc@3_�B��D��5��p	�_ƅ�򢾄|�rR�2"���۞� ����3��e���Ǯ�f��%��u�W��8�R޼���b^D��\� !
�,�g놣>�b�Ω=8�U`��/��#��L*�U5��B�ʖzT�@�@Jḍ@���$y� Y�d4�'�i��N!�j����V̔�����X�pQN��z��w�×�.��$n�R�W+������wz*[)�7^Rc�!��Sk�xP����Y���Ć�a�ʺ���$iw`�1'�'Or�ѺM�ˊ�tZ��7t���k I�h�+� ����UJra��K��]��=�'d�|�Ȏ#�Ke�O���L��;%��q}\L�j�H��ֶ�[��Q�P.W"�>X�/����8\@?����M�|��oo#8$�l��O:���&�,����@���{�L=P��h��Zu�37 ��d4w�^xe
MJ����z����V��K�@��q{�D��d:�#}1$�&Mו�a����訉�OZ��D��aW��%�b�~�(��C�Cu���ޖ�ƛr�T f�)�u����;</]w���t�������ޏ�q�f����LT�~�v�-e�X�K�p��,o����&���SS =>/"�b�M�m ���툹z ��@��7��J�I�Uc���2`�h��r��0R;�6���&�