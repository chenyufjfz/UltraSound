��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ��P�P�I;6��y.�R?* (�B Is.�� �AqQ�s��JV��H��4�b��+w9p���8ң�>��7BHr�3�t�A!���b|���;EܦW�=&�xiC���ցt
�y!�u.e��U�AFx���>��<vѥ4��J�}c5" h`�t�~ʁ�eHev��ִ�X)���W+��0��[M����}�;'�����ŏ�\���������k]��Ŧ�\MVH��������&�����U��ݵ %R�#��
��7������!z�i4Y��4������Z�h��#����G��vѓ�|~�~����^����eD��N�.�k�����*��Mڕ恵���P:#��(�O����d���t�����G�dط"�WЊ���_��K��nVna��ߠ������E��l��y:����z����՝��2i���[� lƝ]�=7T�KG�?��85����k�S!&�"�'|Z9�:���ՙ�:��-]��ҟR����mAH������B\��F�tbӕ*";*>?Av.��yՌ��c�r�9�@�ZR:��}��c؂�e�jF�+�裙m��cX[%,<B�7��>8�U�
�K0q'��r���z�-�mL�0Բ]9�4p�Gt�
��gw�^����h��k,L�=�|\�4ȱ�s�݅os���↴�<�����S0;��_c�Q���r�L�Y����cgX��@ ��;恚�@OjM���gQHW�b_!��i��Z��#9J�k�j�����w�(�Pp������V�XM�z�M�ގ�*;�կ�D�&/h���dE (\��� ,��k����9��ꈴ�Ec��Ԁ��4�+��B'ߤ���tN�!��u�+~�q>���fF���i^�6���I���vi���r�W��P�Ԡ�f�Пr4�a���ݙ��T [O�"#�����Z���?u�?$��n_�tc��x�D�d4;\�S(ϲz�2d2JQ���pߐؑ�g�-��$�ZIφ��>�UK�N���lґ)vt��R��P���D���.	��-����fp;��V+q:Җ��Y��j8��~��&m��-}�_��E�:�es9�=�b��$�74\q�S)�xۧv�6��;�AP��A̻6�H����Xi^�Er�)G�U֦�"33.('�M��`��^�1�7��U,	���WOM)���4n���{���7�ɋ�y��[@�An���"��;;u��AJ��VAS�YQ�ԿV�����I���LZK�Ps"��k�˯؍}�~0A�@OIq"s���e�Zp�3���E����?�x�D��:�O�1�Mڬ����6����2D.�d�OP���Ҍ��ק;g&%Q�$װ����-ӗ�X��������t��R^R}.�b+�?x0�e}$YY�����?# ��n}�f��d��A�6BU^XfK��d�K��꟒<q�(_#�<����a$�j���i\���*��3l����5 &k���lXw �?������;��B������:^�.��R=�D�e{�V���{����J��`���J���91m�D�O�SxȆ��IU�s��%*<�#����o�@�3"3�O�*�Ի����c@4V�TaR�5��9�ԟ��N��\�\�t���I���f�w�1P�1�8Tr�=�[=��Sz�׍�x��͔v>-1������������A�g�3���Tڇ���nC�����9/L��]��X�޿(r�Qx��/L]["/
�m�0�x.���^h��
�t'׸Φy��jL�~(�z9��X��G�j�	o�H��B��,��n(�����U�(��c��W?��y�?+�J+|r��15q�*��=G�[�8�Шk3��F��+�\�1������u���\;��,I�G�\��n�cB
FWX	~`��R�Ϝ�s�<��B��<�<���0#`x���8
���d>���(	��&^n����XJFL�ۨ��E#�u�0���i�^+��fq���2�y}x�M��O���=��9P��^�0^P/�fE��t�r�Ch ��L���σ�tL1�v����&�YZ��s�*�l��]��
P��R�Q�E�	���aN���>deq�ئl% ��H��5[jb�6��	_�wEs�����vv�1s���
�guw:��m��LW����W_̺ˀ�b��+�8�f���W��	Sr���M�����)0;�]�&u�\եx�(Wv)UP>���csނ�4�5h�+���������k�BY��	�}�Q�2�,L0.z�+��ڼ����O9�^_��B�0���WOa�lR�OO�/�Z�5��IԖm�4�����4m�U2�5Xɋ�Tb(��1~����ʇ�eǑ���!�(���b�8$�ϘEg�M�L�O�],���%5n���j��-䋽|?�=�R����8|�5�I���?���-՟���Y�l�|�n��4��6�`z��?.r\���w�Wv���oW#n/���O����'jB����-�M�WGq�=�z����.�$u�����13�F՗��Y�ܮc2l5��N�a�
��n<@���j	!��t20#��"��|J��\vFN߉qc���%�<�e�G��be����lkk�gPD����\D�|Z����XZv��X%��.��&��P�ٺ4J����E�<O�;V���e��h��lu�=	����X]@�ό)��;j�b�`�bhI*� L2�=�]�A���1C�[(Ơ�˪ҧ� Vv�/���Pw����5�@��bcb���Z�A����:~��>u]E�SB����ʈ���%I��V�cL�/��K쟭Ppk�����#k�H�ݐL�8���-���ؿ}��=始��u�z�T��y�W%ڔ*AR��M_��і���}|�J��|��r�a���)�ᰓ}��մ;��� -����r]x?jR����dI ��Y!�C������z��-c���3��ډ�Űb��?)�<�<�/ձ�1@�`xq�Qъ�����R� �m|S�U��rF�����wnrb�+X3�%�����A�N_D,��)�&�/�n�*&�2P���5�����MmZ�yv��!�i�z0��ȴI���������R"�8ʬ���u#����CTob���Dx���Y�����"�]�o�3��h~����p���C.�u�E#���2p�J�1��\)�F;��d�otVҕv�dy����f;I�Y໊�&����(wV�0�	�C����>��+`ͺ�<K��r���P#4���B�P�,mJc�"�_�����Zi~� q)��XI��&�COU9�䶆ι�i��;��B3-�5<�UE �L�S��Fj��������-��/J���i
�\!���&�+�r�Nı�#�HL�� Z� �g5��>��)HЫ��@��r�}��;愓�\3M�ϻG���:��#�S����.��AO�!Z�кi�8����g�I8	�R�q~5�+0m� ��~>E'j$�	j<�&����U��+��} �q�� ��F5'j��	�e�?�\g���Ke�sq�4ۉ��Q�Y�p��%�A����I�-��,��"upp�L�nJ�|ǽxR��~�;��� �D7;
��Iد��'^I�����4b��*#~���u-���Q���;��ؔ��R����6���{��jq��δ�恟��#x����5�����&�R�)c^[�=�`l�p>G��;��M�=|�<^���B2�-?������(q�{a��ݢ�?,�0'�
��i�o�kƂ�|��P�=�" �C��>g���^Yf���a=r��8��l��8��v*<�yh�c��������p�5����U|��Ԝ2fN�p� ���#����;)� V6,�U.�+A�5lr}�ET���tT�T��f�����>;�ya�aE7���#g�*�f�@7L��b��	�ypD�t�­Ë+Axt�Y�´��$ɒ����0��j�=���h
{n�3.G݇,�Ht��P�f�>�����5�Ԇ�]60�'��y�$�6��xfFbZ���Y��"1I��6ss`JG�;!��~>��'G0�:�T���+N{��2d���h�&�~�zCoB��@��x~O�S���x?�S	���DK	�N��BxˮL����`���ǅ�I�w��}á�X����+ �%Һzh4�ވy��X�9R�%��\BF@�`-Ц�Q�?���E��
�vV����8L�A8�)��N&+Wg'"��-%Ǵ��G��|?���t��Q��VyTZ��\�XTM?�j���sp�]A^~���[P��Q3�\Z����������V�O��Np⩇O���Φ,螇��X�4%KR��,dt��_���5=�	�W-�l���C@s8��E���=��/?͛Y�Ze&w�9��ܗQ*�VE&�$�֒ {�����@�~��o���`��hI.ͼ%�)&ʋo��mzE+�3Q���r�}!�w�p�E��9䮬T׼�l�&p�[��Qbi��h��j	[����4X}���z����h��@x���������Q��n���d��*�a:;����;�1�b�Qr��]�/�%'�A��+����6��޵]����� 4
�A�Ep�TX���MB�x�����n����!�	Ч�ݚʂ��4e����(�Q��>���a�>J趿��@6�T���*�SI,��#�u����%:\#�`ѝ͸sD��X2_���y�-����Q��\���C_�SL�?�ګ���z�ˤ��D�bh��Pa��>Vr�\�ۀ�O��S�:N�l���[k��єV~.�-)B���X����{=�[�p�V���*r��ϰ��Hm 4H3�2Y<�%p��V�����}?��W�'l��j�H����zJ��jbg<�����db�'��+h��B�G㣾X��%WWG��7Ne��y�wW�-D_{������)���s�;�|*(G^�Zx6��xU^��߷�4���PՌ@F1���{΄&ʙ�!8�e�!�N�Qrj4�\c3x=�����:K�w�4�/��1`a�hHp�NtT�q��b���滒>S�ݕ�Ȼh�ͣ�`�\8���i��������%9�N���#�В&���y睞`$:���AAJ[��	P[#Wps��н��-(>���?�;��}���ukU�*�:���V/��k�4�Mb�m Aj��!)yځ��Ԧ}W�љ{� ݈��_z�[Ký����z��	ʇfNk�&��[iПFS�k� q�{G.���N�R�O�������L=vu�
��Q�)��W�)Q�<���Ñ�(l�`�,��Bف�1�E���,�U����+늨�V��~��^�m?�7�`覸E�	�)���0K'+#���
]�[���nuIML�d��u.�,�t�T����K�����J��[v�����SL���N��+u!�<E��c
��U�γ5�$�I��o�7/�M�Ԕױ�7�mѷb�K�D}�ʴ�x6ZL����ؕ��������?"�r����ź����{D�h�jg8S�/m��|`������Xj��:��2�6��p3��u4}�Mf"�6-ڿ��]x��u�� &k�L>��_�
26�X<Z�ݍ�j�R,݋	BQws03��ˍ)�e�j�ܹ��jf�����e�KS��>$�_�B((��P�<�󾘍@-\O��S�ѲN=�4�$X���$�4����Zo� ��>��;�Z����8?�L�cWS:A!�}M�%�-'�Ƶ��3Mw`A�����p�1�J�0rt�d8l��3���H����E�"&��,}�K8<G0�4Mzj? ȗ@_ѠnJyrm� � ����78{�z��0���|ϛQ��=r)+o/�(�կ���|M���w"~�T�D���_č�5�=,���6��ayH
7D�+d������T� �J�@�����=��K��c���&���r�/i��p���s;�b�Z���,o�Щ���(��H��T%6@�_�u�@�hN���ȽtI�0׬�#>�&�{㮲�.#A.\�]A�ݱ����2}"�K�u�Z��K��N�^n��&g��:ߪtVQ�I�H�7
�B_#	��Ka��	�뜑�p��*w�A9���ó�ouX	p5�6E+;��
<p·��.X��8o���"�uE���J/z{w���m�<z���;�Lӣ��������i�Σ�M�i㥰קmU��hD������4�F��F]Q�����(�:��=5�E&��:��x�f"�0m<�~�9�1N �O��G�,�Y1�`�K;���Υ��ݷ�,:6W}N�v923=����L�tF�3��(�k�,�˞�t��盯X�2Ls��Y'�ǡ�}4��.��:Z�d=��-4X0|VQ��x��;Yy1��uY*����Ԭ
��*j������-���ⷖf�r$��T�!���6J���׌�/�S����w+*�L�h%h�$}%��EM�Æ+���-�zy��|�*�u�EsWF��ya8�����e�~��4��wc /�O����L�iJ��!�'Ǡg�2�l
�x��g�ӡ���!���]z�8�W�v�.�֛�F`�k��U��Г�5��S82�Ƕ�����#jf�S���h������F+�;�s�V���#wk5N���[�ޗ�*Q g`���UD%
G�X�	�Z���)w��?�q��'���RGC���Om�c07�0��,�H�9+���fR-�E��F�VP�����<�֑��x-� ܩ���"����Gf�&sD�WX�%�"^:����>�A���Z{.���7���6Ƨ�Rx���_?�l�^��X�],�Ca��������6��f�=(�h'D�c��%,�;�G��ۍ
�J�R�T6�;�`A�tt1�3S`��'�1Ij�~���os�GmT�_�sg�X�f�ݟ�_�æB��j���ww[-��Ȏ��TD_�c�E��T��%��.az��]� $�3�����搫���;Q`m�D��gq�f��ٟ��MU`�)��5p��Q�s}�
RN{`5��.��|�f�'���V�����5�ޓ�������$0�ت��0T/Ci�&@*+�"5�_Ye�_����+E��?LWǍ�[�`dF�6�;[w��8�b������^ؙI��g����<��j�������$;��>��;�&�:^��ȭ��EC��P�6k���w�F����W��$}����Ӝ��᳝Vg��a�|z(�`߃X��l���op.M�qc5I�y��4�nO!�|�+�5��܆��4|��k��WV���{2!�Z��ë�!y���0+�z~�-�~�� �U؟Ȼi��=� ��[�w�Q<4{�����rz��}9+� M����?H=]MX̢��$d��$���(���Z	i��Qe��\��8(��0̏�>�_��@�Qk�iF�|�ްj,o ��;&�Q��C�GQ2�V�_FV0ʵ��6$y��1�n�'��Y̓�g���T�)�~O�Od��@'&˞�1�bx�^�� �T��t8W����
<in��K�m%���4)��Hrsce����-�u͵���vW����,�`��@H0�Q��5x$h�z^(\�`���ϥ3����&����Vы��0�i�B��o�E:��J������t���I�7�2S�,�B�y@2Z댤yE�f�=O߿���tz[���OZ���t�wݳ�.�3���5�D �E1�E��l�⫖
��3��Ӏ��iM�)�H�_'��f�����{J5������F,z�(��oֺ!Ki��|x���k�\M���ٚL&��Py�����@Xv;�膦�	�p��5#ZK�r��IT���ә�~�fB6Or�\�|��K�DͲ��T�]�<�,�k|{`�ʗn����t'��鬂��T��3�tr����z
����,«0���^�H>_){�4#�{��@4�W��!u��=�"ĢD�KlI0�}힡D4m� �7���V,o�Kz�������2m'����R=9ȶ3f�l�fi(����\jP����%������X�
�n����OH�`z3�5���t:rE�}Z�,�]|�'�Sh�;'�aC��O�7�5�۞��j+1(��u������gM��*�yU�dl�N��f�����1s�vz#��Q�`b���	J��y�Y���^{�Lu�����j<mY�)����3�H�i
[�n:37�0��0�ai�7���.,��s���k�RhED�jҾ\���W�uZ�6�'��n���$�s�Mm�ſl�n�����'v����_�i��>3[AX[��eA�ګQ����=/�[���٪Ϡ�W���+-+jMs�˪nc�4��aI��N���w��u`�N3 `�o;	��Π�c�:�Yr9�	�7���y��0�-���Y�h?�t��7QKS�J�jv]�j�4��Eo2*��2s@�I�������U�[G���Jw���\�3uE�8f���IHb�MZ⌰7�Kt�g�L`��A�}�_�jn�*0�}O�t<B����U��3�s��1ek�+@�%`܆"�?\����*d���;k&��O����i�g�I42�Ŭ�#��9��0 �<�����u�\_K2������Ԓ�'nΞHr�?x_�?S��i��`lMc�q���ߒD�H��/P���E�Xx�����,����D/ba��iM7�e,��+��@�h��;�G��i������@.����
|;�My��]� I�ݜݴ�1zgÍ���n��GBv�V�i! S]�%0�N��j^���|��#:-�w�i�ҦC���tA�Wj�M@�a�h��0������d�����y1qdb�W�]KG��|�)��oA�����݋6����{2!��V����p�GE1�m@xr?Č��GTIQ��Յ����y�@��z\p�$��>�*�_Te��J��V#EKY�Oz9شKXù�.�!}]q*j�؁��D,�!��'�.��f�k�>^U�~V���}o �Yٰ�^	��ce�C��-&�$�8��ζ����bes�	�t.��HV���@eril�`���|a`���>1�x&��.WSJ� ��������C��y6U�1���SCx8۫�nݹ��._��s���x2���J�q��/����?��tbfY�7|�8�W�v��`p����P�hz���a�U�뒟��C��'(|\>T�a�V.�Z�dw[W�m�)��O�蜱]�~T��3ɪ\
� +�t> EAw`Ԏ�]. ��J%�8;9u۹��=�`qD��,���k�T�8�b��PH��D��A���lG���D�*�bCα\o���o4�$��y��ߩk��8o�e�掉�TE�_��o�m���Y{�K�y�� 4�
��N��n.SS��������bk�Z��C��K�<�K+��Z_��]�J�4�տJU)16����ND���ol{�f�r�ـ�0�1��#���&{��2J@���D�]�5>�������F$�K£	fx��-U4Z��}��X�A�`���X�Vq�����Y�N�6�|
9ow��K	
���� ��1~r�b�nC���s�ɑ [�*�)@����f_y�j�v�|��Ӕo�O(�x�\�-+��
�?既U�4%��.V�Br��W��xc�҅�������;G�}-&�]��t3y��[ Ă ɞ
R䪓�"�� G6l@�e�`P2-
	��82�ꡧy �1ˎձ��lxsH�v9�'K�IrE���w!^T4�; 5fbw<�d?� 1������れ�������z5@�^t�<�qu���6�3L��Ov�C��B]c3X�p�;L�q-���9�EN-*0咙.��<ΰ�'�H���2��k�����=��1��"��n�J O�yQ�V��-NjJc\����F+im�~)�'���v�a�$!�`!JԤ��~v؋}Yִ{d�3�B��N��� �"˵�?�Ĩ]3J��b��R�ViE�\��7Üh��FJ���� �<�1J�v�}�CR��y^�S'��VB�"0�D]�\qī�v4��x�f��+f��)!�Ղ�e�B]lհ�%Y4%]l#G���f�M� ������D�m�mϟ�Ծ�Ra�4X��g��ĉ��Ѵ�wr�^:���
`0*�g��:S�6���6I*?�e�����D�a�TK�^�a���y��'2y���W^^��EA��hyWK1e���� 4�<��5=趈@4Y�?�]�1�e�,�
x�#��R�Y?�$zNm$>��2S��\��i3D�;&�{������_έ&;�^����޳���K��͌�t
���( P�Y8�D)ͭ�/X�Nh����w�� ,���#�!lQJ~���:J��=�Ύ��"�o3-�N��Y}+�Ǌ���T�we��D��y�a����*Y1�U�e���.L�N��=�^�b|���yad����F�#S_	������[��HT��%�W���؞'��g�yq�vh|��9��r����YnE.�S>h�mcA�)���uc P�p��m��=q�1k���V�P1��iX&~	l7DU-��f4}C%�����gX�p�׶y�*��{`GDG�J�kv��pW�V.?�!n��.�M��#7�8���%NN�$�s��;;���}��H	IL�t�����D��@��b��}D��d��w�*�}����?(��yޗG�"��oؖ��|��y� ���S=\�"DE�~�"暉\��SW>$�;��>�1�U~0Ѓc�D[���Rb�6#S�@�p��R�y�ld������af[e\1S��֍^�젗-�u�r��-�m�Ͱ����^W�J;@��d3~�fE_O~ۚ8��2lf�(�B��ü��T�qk��r�Ⱦ�SFe���S����j�^$|����YEv�(���uC�=C�@�L�S�'�������@9kg�W�+dV>�3�͗6�#�Aa��H�Xe���>��!��3�L��jI�gZ���ׄ����c�E^{�=`��ӝ��k���$��G�	�Jf�u�>��}(�bڠ`~�{4ε�W��s��܎�=����%R~y���2��ɜ�`u�Q0�_~~���z6fB<% �?�=��W