��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�
���B�+,���O�t9�������-yJ��N���Z��?��c���kU��!�j�#�JD*�������R?�uƀѽnlH��߮ؼ�����3��G�� ������C��w�6��*ʺ��?�1��+��C����챇�LII�{>��g��<��9���%�~��ݫ���v����J�m/���{� t�7��pI��3s��P��.��p��%H�x�>}Pn%���k���J�u���&�f�QΈ�9�.T�8��%�z]�v˗���'�/7c��b�H9��A:v	o`�o��RA��O��������'��K50�?�O�?�]��l��:X �}���s����z������}|=�a�8 �rNvg��o6�k5?�FVe	/)�疳%uwVJ���䓄����r�=l�w���V"�����ca�����v�����a������!,��hy�ڞ�+B��}���]���̆�6���?�W��y4կ�^��iU9 �l�q6�u�Z$6����㙂g���67�m�4��=���RቋU�zhW>4�H���
G�C|�l���(j�]�Q0)V�1.�?��;��A[�䡏EĹ8�ƙ/:VZm����,�(J6!F�T�ua3��Q��V&�9�I�Q���|���N��o��:> Bm��UO���
oUӰi���4��:��I��ˬ��ߴ��$sx���j,��z��N:�p��W_o�s<�'�Ԡ����Cb@[�X�6o��V�%���"�Ǯ��80\�}��U���Z��Y��N5,I:yW��~G ��Â��-�|�q����d�� 3��A�/���M�Ȥ�t�mG�@i�	�2l����A�2��8�"ө*��vL-]rQ�4D��Ȱk�:�ZK�5r�W�"pc�`xaKb�(�ӿd���D_�U��ز 8�Z�+��W��T���Aunc��)ڛ�|���W*}�D/�&�ш�y��*d+؂���i�NjJ��;��c`�G.d}-K�T���q2��o1ZHњlX~d�:6�3�)п��՗�e� ���;C�=h��:y�;��K��dĝ�n�	��rǭ�B=+����&��v4�RxH㉢�(�ّ4�WpDS�����`ʭm���A�JU:���f7�����x6�77�']�������&�/�ʥν\�ߜDun �t����B5�:��P����-��Bf�.ܪ�n,�����n��=b����N$BY=`wh��l-i@�.�g"B�'^\p���)�B��L�aa�$\��ʢ|�S��VW	�؍:�W�	F�{.�c��K���_��Al�����U�☦v0O��v(ɑ�jЯ(H{�e]��2pu)�R�é�LH�k�+߰�poB��i�u+ yü�M�5����E'�5b>�s��k-Z(�c�|<��h���4�dȕ�V��=�;&T���v��P;����W�-�n��hƮڨ:���7O�e�;<��۾�ٴK�"f0`'Ġ��D�J�ĸ��{>RbEvs:���f\�'�5�-$��)�^�h��=�T~Ǚ��⫣�o2\�c�����mq�L;r�je��A�k|X-�8,K}A"�����ޙ��Oj�^����)C��c��1�u��up�с6�M&�Ȗ��EID[X���z�(\$< V:�82j)�* ���N�V
�𲉟>�c����4��b�.~E���2e[�:n�Q�Zx�o�z[�'ܗ�Ъ��������>�.���48������o��~G��hR���)��ٶ*d.Q2&}P8�4/���L�0@��U�k�?�HN2N0��q����*Ac���6G��@;願Na�	�`������HcB�N,|K�V�%O�g�u�5�$�0�	�B��eƺ�H�.e��;�.�HM5_k$�Z���&/{��~��J������6Ї+����B`4�
���ڠ����U9B����^���n��w��m�;������`\�,�H�m����ޣ��A����MT;yă9����& ��t��?3ɔ�`�P{����,����b�}8�6,��BR�ip��x�]d���sJ/���D,�48A��qh����ӁO���oA�J0�E��Y#e9�*KL'O��H�D�(��	�F�`nx%�Ϗ�d �����ȶ"�9��,�k��>�g�TC?�$!���ә�nc��t���K�k�3�7g%��[P�'��t�Ȁ!6(R���F�𥳦� �<DC��|i����(=^,V�e5��'X��W(&�n�^�Ն�k��Ra_*i_]�(�?݉ ^�ՍoA���;-x]b������}Cٻ��#���:o�hݶ��j?j:�&�S6�/:h:G�X��Q8�F�����..�\J[��3�#�f�X2~@M���@��+�f��h?Z���O=br�p�,�qySC��T̃��$̚h�����a?&|C8FXA��Qv��f��|��I��+�����긔y�����ֈ����Ɲ����v!n`�۩8di<b���D�����|��E�U�l�)�iFm��i�e�/�L���վ|���7������	CIѦzֵ#^f:���w·�[$;2��d^�#��3���A�u�D���r'e��
��d�}_n�"����&��ܺ�s5٩�`k1�1��2���I�^&p#p����@�֎E��9�j�F.�����P���0Sp��NU�zW|�&��ػf�(nN$#;Q�n�EE�l-�m6
���$�wM�y��=u��ֱHC�MS��<��)֟���]�@�����-��|X��񖯝H�k��-�I���@T�ZA��ŴO��n��Ţ��v1 �o���KW�Vqp�>2p�~g����6v<���~�q����o�kmׂZ�j�]�g�!,?;A�Ö�f5�P�rᎊt�]f����u� W��C<٥�	"y�^����~�g/NVGGq�[��-�F�t�4gtG���g	vx���G0-���pEpp�O,�F��o��2�/��V��B\�3�"k�B\a��c���x��Z�L�M��C�kČr�?�8R賽�t�-�ܟ����p��Bӻb�vL�<չf)"�j���⛄@�:�&�ߚ��9#8�!�1��T�Z�JO:�3:-�G�mBV���|�[���d%-~&G�B�����\e���M����wE����k�TE���
���jM
��Dͥ�p���K�����Ⱦ:�~�r�进���%IU��I/��̸��������^��V9qy?/���.�������:�e��`��q�v�劉�Z.�a���ܬ�;�|u}��M�z��Q���u �[�A�����X��f?����Gv��ݲ��D�w�4.�Wn5[�1I9W�[���Pa�ᇰl�6~qRĖV�L����_V62��WN��IS/3Ɨ��(90���S'����E���횚���\},�f6�b�jK�͈�$#���)�K?���i��|ۤ��������稧K�����]QR�����1#�Ig@���OR_����aC��t�ɽT;&��E��=����t������͍n�t=�˳�^�(�1�y.���䅰�v=��7��*![;�3��C�.`���ݴ6�^J=�1�������4������]�9)��%%�֠��,<'�_��A�鵷�d4�Q���z'<���	��B<�M�y���P�`��5D��3�&��Hù""��0z�u?�Be0T��#���~r�p�R��j�e�XO��-Bئ9�!�/��6��k�-�T��\M��Q!�, �C6Ŧ�R�3�t��(CJ�e7�kRdo1��f_$QXN�R���H�f��zB�"J���g��31�0?.�2m(k<م�fu�X���z�p��A��AM���k���u���y�2��?I�,�ХfjT��D�)��&��g�% ��U��Y�����9�����|�?���˪]{e��7%���ђF^�`GF�'������-��Ӛ�%�ɹ��]׵_�{����L2�[��ԦNqg>֣x �3
�2ys�9��Nf�X��뢢l'>s,I^)䫎��'.�����8��:DE�َ)IO�]s�vI�0<EZ$^��4e���o��«8	m�	��� z�y�Qjܔ$��e�+��>�����8����!t�Y�Dn��l)��I��;w;���pm-���4������� ���b�.�}�����9��&^}��A"�7GE1C��J��y�@�h�G�H]����B~:�ud���8��i���oY�,"�n[���g�� ��\�;���+�-�S�L���UP��F1�FЇK'�W]�S�X�jV����j����i�=Rց��N��4���@��F5(�Q5@-�=�R٩?�KJ�<�jWZ�N���H�x���'~�^�ɶasBO���^-7�~��/�ɂi�F�vpW����lU:];��ĕ�
b� K���l��n��j��-TG�8æОQ��/�=�!#����mi.#��a���?it1�P,�n�		�Q��0�����+,R�X����(?�x^������]�V	vE�������7\N��?FG>8WQ_�L�v�����E���u�L������铌�[Ay�<�1�G��	��K?.�Gm���<y��Y�r̜ҥ���;lS4����Ty�_~�kZh&��D2��/")�x�c���p0� Ȩ$���P&�9�KX:KJ����f����Y��:���yL�+Y����s���D�S��oĄ����S!� 
�%��j�~�׿�� phmp�Ƃ0�$&*Hq�
�{]k&3��(��1�����X���4Q3�T=g�;�!�>x���i��h��s�L����i�3_�E��h�!�U����L��/��@1m<� ́c<QB�}��Į=��#������	�~�1:#��oNס��]�GN)�K�w�M��aA�DT���g�����6���=����4�:�����?:�ʂh#���)��3�S�$e�}sda`���p+��#�}_�$�0'�j�6m�o�}�iJ{�X� ~��C��&���ֳ�{��(�_.��f�f����s���Wl����'�IvKQ���!(��%.�vi$J� �E�ڀ[��`IWE9ķ>��G9�yM�W|*���N>�ꑟQ4�i�eշ�<�$_R��
v�$������&�2F��RG�u�2�&��C������zU�O��tE�t?&���Fp�������H�}0A�h|r6eW&
����(��r��l��4��[W�%"v��|�M���4ek��Y�n7H&��q�|<5Y���©]ۚ\h�ʓV:!��9l��K���R ������'{��j���l����$�@���R�>���P��J~�6�a����m
���x&����]��Ǹ�;.�B*׀ou�|~��� �]�=�^8w�W�գ���u1�tPƗ}G}��C2.Nss]k�DL�0
{,Z���hM6]�u�!9�S�ą�8w��v�p�DYU<'�P��qH�3������`ᆷr�D3�V<��V.׊��Mm�{�O+��� BsD�|�,FL��[r �g�c('�44(4�M�X]4_����Դ����A�#�6f7��g.�4���L�[�v�X#G�
�@w_jX�U����I����r=9�?�>�
����2nz>���/�Y�w}�X�I����I���NV-/kVb&f��s�s�i�7Ӣ��4�m*��������T��)�-Վ�����Z�ձ5���*Q	�E�-���3|\��UX��Wf-L�0i��������+*���Sr�&�s cQ���zX��D�I们�p�{t��RV���t�\��Җ;c(���p���?V�;>����C�9���l+���	��kq�&���,�w{���i:��8T�P'v?�cUbu|����1҃X�=j��G��m���
W�R�"�&ͅڋ]�w�	iZ�ݪ}�F�͸�
��{C��X�X�U(�Hn��[$�M�a�E'�e�����y�]���a3��w�H`6�-ό���`U�o���Fw�yl�Y�O	p.��`��/�Αz�`�Y9������ش�����ȁ�A��o�����j�V=����R.fA��`�r�� w�*�#V/\t<t }��U�?h�q'�$�x�"x������Y��xAp�$d6��f��'�?0�0�] �%��M�N�Y��8�9B�r��v�E^8�%u֝t�5hS���0Y��l�Gqn���(�H:��\�F�����0`�[d�<)�d41��q+I|؊�#������V� �L~
T_4��)eX��:���
��Q��t˱����9D��-?�X4Q;N\Ǌ��rĹ9$�xu�HLmP�A}�A�y�Lb����#��O������D��R&$�+�'�V=MYk`U�Q��^�9azq(�V?e�k�ϓ�������j��G�v$F�-~�����SpD����lMk��F>�v��[�J1f����v"�4����4H>�%��I��������3u6!B��Y�Q3�:��(��g�ӑc ���¼�!�0�K����~�@�PϽρ��J¤���\.�a��~h�`,l�� ��0�(���쪫�>���L���jH&`��@��hd�cWi�Y��j �Od���n�vO��+���dk�uO���D�u�1'N������_�7�b�
:~����
��v��u6/8=�.Etk�P"
,6?`���q�ܖ�}5����HAU1c@��9q3hSg���*�M�XpS�`�ꪗ���B���N����g�����q42?T��s�g�E"����?���k��q�"���&@!^��_U�w=�t�IM.�۶cD8WPK8��I���"����&�_��SfP."C��(���N��5���8���{zL@��4��.����ؐ~ÿj��s9�dw%b�&=`��� ��%�_�b��c�4��zz��C���nd/s_���U��9��&��+�� 2o�����>Z�P�&#7A	<��\����Xj��2�;4@�MA����Ui��F� �(/�!D4�efإv����
F�o��t�)�H��ն��F�~C��Z	�B"�٭�u��������y��fJ|��e<�ɦHs%�{d}틵z��_"�Y�jv�,�l�1�ަ���'=ۋ�Z��[jx��o�+��D̸��/����qKS:Α�?����{�����=�%��ѱΤ2^'a�D�<pXk#��)�)ch&'!4��܂d<�&5 ��oDW��=e�Sɫ&����&uS��}?Ŷ�Lo�N�2o��\?;��u���9A����/d����b�Z�;��IY�<e��O#Ag�C%�(�
�A�T��.�/��R��4�jn*r��K���X��z��V��=!g}�p��)#��A�$"�P�I��Xp�1�+�&�����pr;Y��C3G
����r߫Ì*��*n��:�0��[�m��,�k-��l�[J���>�?b�4O��wC��	�,��O����m�c�5%u� QX2��n��A�!���iyн�\y�,���s�@w�v�B]>=A�0�'>�!�T���?�y0�N�F�����Y/���j�_r��0���O|	�f�͑O�
��I��eף�3Y([bu�<���|p�%9��p@���j�(��`�D���e�q��������:���ó��:��[�cz]䲂�U4a`_�oq�s�b\�z�+�&�(D#?R/P����?�
Q^�z�y��E���xF�r��*\�z��-���"��]L���|=Ň ������/(��T4�O���p�M�܇M�@��Kl���F�M�^Rf����Ys���ߟ�R�.�I�,@� 2M: �ݓ#���ԟ&by2 ���<����Հ�e{C3Q�Ѓ�"|�r���|�#Gd$Wf&���~Ɩf�p�q��-ư`�'K�&�?�T��h/]�h������w[V���FL�h�ZV�����|.�h�imڒI�!�3\3x�w���t�  9�)aT;�	!K�и�2?jGp��¤g��=T}�D&Ǚ��h�?1�����%����S��~�	�t�pLC�״p�W���Kio��X;'���� ����R�t��\�w5|�O�
���̤S���\Ώ*�6Ubϳ�>�5YX�-�V�(�T��}I�<+�V�7R�^��M(�!�;��3
��mpz�V�@��$�|�Q�/�,x���*r��W:��B�����Ox����Y�
:���.�3���"KP�i�K��4�����(FVT�I�%��� ��)Hb��Np�y�X��]@9o�]��\�@׵�r�LN$Jʇ�+��h�:��b�Hp��R_�Li5�|�K����ԳH������=��_�d�&*A�ukb�w�z�<������?ec���r��`v�!Y�� {����뉉!�.ᐒ�)m���4����SԀ'p�0I�;��P�u��}���1D94���4BQj��Y�Ӌ��:<�cdd��Â��.�R�i����x1j����{��I~�'���b�"H�i��x�V�	�x3�guI�vdJ#�F f,_��ۊZ
����5�zA���)aGM��wn��O���bx����[�c�ӈ`��_#~[?��^+s��s�_���[�H�k} �8"�`�)*�Q�� u��H�D\�N�y�%�
��W����27�6 E�#
�6d�s�
 ��]ؗ���,%�)O����4�w�}��}�7�h~4�*�마�b�uj!7A"\�n������c:��2#nE#-p�k��@�豻a��u�n�(U!|�Si�[^��xf�"=���5�{,D�[v�u[Dғs����+3���Kټ�PZT����Q�����VO�F���L��3���X(q��]��E|W���q�˱A��,p�G�qW
��n {�Ƈ껰�$z&~���������͂>�MU��k���U����~( ���"}�:��t�C��ň���&��Hgý�(]�C?<\�	�V��B=�;v0��+rؕ�w��T��y��k�&�M��A�~�r���̌���m��r�V�2zrڙ�b��v?Qd�I�.������ȷ~�����sC�o��gYT
�-�]�(��4u��Q�:�Ni��� s(��|���Mw���d�%�K0����q���b��B7y��ۺo��Mj�Ei��M�.��v)S|<r!��q��y��->�׸A��z�!�W��q٭�PP!vZNWo�Ǎ~I=���8�������7�]���QZ�=Mo�%8
�s�*�Ά��%"g�{(����uK�kݲ;�]��>�P`����9�������G��i
`ʞX����΄H�R�_�,}X��Yާtd�n��]']���^ oST�W;����D��-�"+����/�|���Ån"�p��s��IW�Ą�%���M�&	���	q���������0�I�J���zZ�����a �.�%�ͯv���	I�{C:�\���#b�u�^HK�j}  �xs�,A����SF�\���$��|�lٚOD�vp�3�ר���MG�3\~sO�?k�Y�&8�4Ib")�+����Jl��:+�Q�$���&�~Dp���u,�~_-�|Ee���K��`�A/!B)�����I˰�K����&F�A�S���%xy.iq�����~��.;|A��l�?�2ˋ!��Ym�G��%؀]L���|��j�u������g4H*����o�ċ*������sΎ��*����#,���D�`��.���� ��Ѥu9<5)п�2/*�hI�׹x������+J&@V �ҍ��+?Ǹۊ@"�Q�/0,m���u�h,��;W7<T8C�HP��9^G�=vC:3^���S�O��	��d�&�N��e�{�.w�A��O���'�'���{'̶��I�;0�H`Ρ����6��u-
�o��mW72��Rs�h�y����Ǔfw_�Pa�^u"��B�zw+�-9¹ʟ@6��8)���dա�`�����Xc��yJ��.���6P����#�؜��/��b�d&^K2W���P�Ȥ�ٸKK����˳rk�yz*�_�iJCH�K������������g�ӧH��� rV�75�A��';�^��#�.��@`�o3+NȊV��2<Yo�#��A��x��ʦ�J�p�>�	����QquQv"]N$g*]Vk�V����=�0P�����P5�\s�v��U�k9�y�L���ı����Q��Tz]�P�h\2�\x%��ֳZK��[�����v�v��Z8@�Tn��G�J({O��#T����:Ӑ�b�낊U)+uS��pP�ׁ�H�Mȁ8X�	4�J�ky[��s�8?�����t���6�	)����lq�a���	:h�Y�uSc��yК�h-Ka�.����Hgyi���>�������<w�9yX�S�hOq"��L�x#$o;�?[�΅A]�L��l[�PAF����Gu�5j;�\a���S�Ѓ 2��@�/Z�H�[}`�B#��Y-6z�j�k��e�p�=�.gy��{p2p�v	�\?�.ӻ�יW(�Ű�T�K��L���a��L�2����f�~P;G�O3�z�$�������7b���.�{��S���ńh��j��Q$b�MLB��V�ҥ��'��2w�󡘟��/���d&Q���f>�;��T��/������h``�������uXm1�+�;nC�\/�lu��U��������������2���#���%�:J�sFc�V;5l�i��oM��A�\��Di�k̋m���tW^mH�IA�tf�TZ�뀄A��p'�as�Ep0ق�0h�4
��b����$4��hlܡ-hb:���:�4��4��Q��w�F1朢(�tP��CG_H0�/ K�c7�kes�qx[a��|��s/�S�L#Ly����4?�u�V/�|���d�Y]�K�K՞e�����-h}�����V�U���tn�Q�P�Sd��mZ��F�B�T���T�7�Ґ����.��gF:W�6����'"`��=�X�S�����
�!̲�M��HR�VUu�~3�Ymw�X�������*_����)�E�| �Hߙ�lz�����n�X>�48�m��3Ϸ+ZG�UR� j�ۋ�����z�_��E���$
�w�o4)�㸜~&c��i����VX*�L�z���=G�=�	��jKߨ%_�v����u^:f�DS�e`m�ً�d��횺����z������[�j�M��(����m@�!�E�ɫf�xZR��~�È7��va���P�i'l��os�
:���y�J������@���S�L��DZ��5Ʈ�BM[ה2�فXw�b������6�]��e}�8��w1�S��/H�WL|�
N�t"Tbޥ��_$��㧳1�M)�����I-�ثV�{�zx �Z�h��4�mVa9�C�\{��q�SY�r�]�I>kX��!�}2л�J�-���!��~��g��a1�x]k�?.��z�3�� �h��{� =�,8��toi�Q���ob�-"s?f�fyb���tx�O��H�[b*l\��v�o����B�uk����٨���rq���m�;�����A�?���)ff�ip-w�fq�W��3�A��I���;��d�����5�����_���;�Z�1 _�"��Y,�r�b��9�����y�.c�^��l$�c�ôշ�?���22��d맙x�a�c��9�������H�;VLњǡ쑌m���"h������6FxB���$���l ��go:�+8��?i���P6��!	��Q	ܒ���wΛ�\�n!I�@UM?�9	
��ɶE􎐾��z�&�37��9����7�Ю���ȏDJ&�ܻ����jɢ�1*����\�h���NP�:���2������� 桕�0Ѻ�h� 8U(97	t7�Ah�dv�Ĉ�;q�m��=�ԍ���Ч�k�>wӗ�=a��(z�e``�]7�"đ;0�CV�+Fȍ6�x��z�Y=��Q��P�6F)!

���i����K���л����&��)7���A('˸��@�t]���T�����1GW�¸o�8�C�JZ?��D|����r��}b�q>���㼔�\<.�Ջ��ϭ�h�k5��4��-�i��g��
�� )VR�F[��'� |0�)�k
ņ����Qڊ[ذa|j�7Ɨ���]xt�9����om�I��'�S�F£Q��=t��ۼ�[�F��(ć���}�����uCґ�,�����&��cXg8��pgӇ���#q��y��T%��SЮ��6�f5�O�SH�C^FE��~�t�o�Y�9 �?T�ZE��,$���˹ɐ�I6�@��Zs��\w���r]�����< �}@���_DW���I�A���x��^�z�.��R���ؔ��U��$&�C�瞛!oN��~��4�.��d���W�g<R���]��`�?���7���-�#���I-n�d�t�璻� T�YE�X��>��=����X�ҝ'�$a�K��|zE#բ��!�0�j:(r���Z���g�h���b�l�������u��F����Z�y��3 e��yr�`/Y-w�\���Tʰ&7f���N����2v�$��� ���M*���i?D��XTGv��3�:�f<\Nߘ����}�FM^*���Ir� ��nWY�8�&]|۪R��F�F���ȵ��O߈�,l$���֎�9h��*N{��c���-.�P�����B�%����~��n<��LeWᢕz�2\VF.�'�)bm}ǉ��4`��h����*��rx�(R#]�D���ɯe�P~i��u����yH�\�S7��O����e���P.�5`��[?�/�V���E���g6]��\8�ު�5L���,-��g/��z�O��UIsE�M^"8��3Wt�ֈ���z���=%*|�BZ��~�A���	J�]�fo��5��3��❤�'�q��qH6�%��l�֕��d�&+ə�ϡ�oTN��7��������Q`�bzy�F�Wvl-wD��V[�%��w�=��>="���v����cKܸ��C������f��@���},u��£�W�qВ�ˡQe�.I��P�]t5YC�c'$��`�3����[���r
����]5vߋ:�G�Ii�Ȣ�����󟻳���7p��g��q�h����
��|�*��W�7��:$�Gi1nQY�|������W!��b�ytD���*'�U� Q��^�wf��;E� �������{J��ߑ�.�jyw�Req�;P���'\��E��a���>���+����2��)o�T�]��9����w�H��a ^���	y-�?�����9?��Q��ɓ/ (X�?Qv�&ޞSB�R>��b��9��vz�Ͱ��"��H�|�Z��Z���'uh419K���#�{������%!.�Jh�63-����Tg#5�7�MgtX<�)*����Γ%�\�pTЎ��B�'yq/�t�Vvn�G��l�0'�״����D[�#�]��NΨ$M?�����o��N۷�N}?$�+d����/�_*�%5x����Cش͹*'v�%�]A��&�����-p�2���Ƨ�W��oH������ԝ|k�p:�u:347v��$.R�{(�7��a���C8?NP<"�ag��a�Y�?
賎E�U��}���A3�t�=J>�{?�%����w�}�a+v_c����>s0�D8����8�I7F+��;��(�0��3�df��L3����9�T���!x�X3�@I�V��< �	�y�^��1�<�IG��(Al5����x�9gz�HW���-�Gl���s\~�5��H�/��x����7���D���fc[�>*�=9��%�q:��H�,�_(�Z�A��w���>��z܀ǵ��F �Ұ�%>��������A�"��(=^�v��k����_�� H� �9f��f�2ȋ~G�u�0Q�&9i�����b��_���A��#��;���N�I$�)�o�G
�78���?�5��"��U��+�k\�8����_�=�����W����tpEn"E�kCc8�����W�Ubы������燌]B)�����w��<q��J�(���~M׊x���.�S�l�:ߎ4��nI]��~�����(�+�\;�&����r���i=��5�~#P$�2�I`�R��$v��!	sz����3�!�	d��d��@_D�k��qX��V�"?6Ct��bR�ɍ6��&P��/���ŕ1�z���=�ߑ���k���Z����`�ʽ5!d/8��	t�
<����k�N<z#a��Ƕ@#�6����y�r���T㍚������_�i�D4}q�1Hg.�����a���N]�4�ƋJ��o�͍������w�p�.�B&M�NvD[0c��	<G�,��h��G3�
�Pv�ԬFK`�Ǭ���O��?u��}�W[xOA��8��*]���]��.o��F#������y�=N��- 1��]�K����� �]
�c)U�*��������c��^� )H�;�T��_� NmJ��������
F�$��S�.X_X7ի�˂^q]5hw�U(�ν�r�Wӈ����-��M��<�oG��K�9���(��~��r�$�����ޗ�huÑ��<rE�][a,ˉN���>��^�?���~�4�]���� .tٜ�u�#��N��SXz���瀬
�ӕܷ+�f4rmU}ꡚ R����0g& Yǖܱ��f��4ᡰRˎ�*޻Y��b���7D���mu�m��mc�7�h$)~��9䋶t���E�6н�����t�V��>�<�
�H�躘�o�aPl�g��'O�V�~n��c ��t�1�P��˜��B�Oe4y���G�}Q�}.zFM�������o�:��VPp1�t8�H���?n�p|���OK�H~�$���,�J��M�tކT�O5u�:�`���̵J��"�.���͔N
����7F�!9�}\��e�O�aeB��rx��H�A�0u�+ޖ�^hLd�d_�q��e@Z5�!� lW�?J���\9
��j�_���K�av��Xf��"�Dk�Y��(:��j�p.�ޑ��A�HJ�9w���T�Y�U�y���=��,���Ӄ�V�f��P�F�M��͈���i��r�4l�Y���P���Ж_\/H�r)�B<��/Y��Oւ� nb��~��z~KS��p �?��r30	�4�Ǹb1��N�_Ɏ���%��MګH?�?�|[Jئ�`ԫ�
zc�����Aʽ�1��Q��/�{yiV������;$�B��K>��(�W{Pl#��-�D�q\���9�/���*��h���l���[ցwU�C���ߍb�`9��xy�JY"? g�s���Q ���p���)t�#�Z��'� @#��i+]�V�ǩE@1lT��7dT�sض���U-�#�Y�Wk��_c���n�H���.T��c�N��W�`�T�Ihd�aSt���`���^1`��L8�CC�/�N������n �����KI��E~<NͅV�r���8���y�H=��Y��V�;�<�5U��f[��5�C��-qr���2����둣t�*��yp�A��FY�q��]P2,y�a��ͿWϠJ���Kv���D\F���ԫ��)F��2�҅��a�+��8K�~��Y�T��V#����vP�ѷ�+�"e��s��ϑm8���
b�M��Ձ&v%1O��2�(�S� ��PX�<Z�J����ߐ+?�`e���a�~�B�����X=�pE�{���BC�^��Z!Zh�	mtV�ʜ �1C�(���2o��P�!��0�W���'� e����zysi�GW�37|Z=쳂���9���� ]|sC�ba��-a��M���Y���mO�Z��O�uc7�+-�O����l>�oZ��5ti?������oE��0p�n=Z�<����� bx���ݶz�U����2P��-i�1�z!��w'0'@'���g�{�S��Ս�������dycRZ�P��|�Ӯ���w�QduZPfT&D��0�>�UFZ�p��>1]M�=`A����iڊ�ەL$16���wM�$�ƕ*�V�5�Ҿ"��5:���Ir �=��K�Ӧ�O<�PQ�|e��߮!�[G@% {����z�y�@��^kr}u�t5�k�y���&�\#I�T��
�x�s�+pHШ�+#e��m��baP���e]kmƹ��_88j+�q����:u}ێ��c�Wj�uA�;C+�?F�F�G��/v{)W����60jr���-�,I�cB��M�~ʻ���`m��0�����K��rZB��R�t����I�x�IԱC��D�x�F��ڛq��-�F 2���e��H�>��i�#�;K��#r���������0!xٝ���ϔK�G�����oϼr�hV�7���P^5!��8�؊�O����b4x�&ǚ!��T^V,�p8�a��Xw�mh�k�o~ܪ�@��>�M��B�=�
�F���WR��_�O��ΌU��U��y��?��a��	��"���qŅ��yY���.fؾ���u�~1ہx= ��jS�&&���A����֛��p�6���7�����4��'S�J�4�	��?��ӷ�p�Y�%%8���|��]u�ρ���ѷ��9�`�y�;�[�u�.I���p�V_�~��%��KY���Ue7XAl��j1V}a��L�#����_mL�����Zc#��w��H�kMS����a�(}H@�������Y�J��CѐU��P���JTU06An�FX+%Ɩ���~�2��&�t�/�OS�\�	�2uxI#��k&ȭͳ��Q��iV�^_�6���6q�OL�@T�bPw �]Tc�{�����c��֊���h�MIH���F2|��M�,���G�2Hey�����A)\D�����{1MLw
��@���qu=��yɤ��559�?�/	mL�R�.��:�P/y���G����Xh$�aR��7AQ�f��bO����j�7>��ۈo�sE���s\��J���n(q����(�A���f�D���"Z�����Y������Lwu��A7�hR�!i�����Т"7��E#�������ڣWj�FԻ�9�/��T��t�'f���D�����msR��϶d�5LEE�����h���	�,`?�@p`���<�påt�r���ƒ(�@����mr���r\����h�Q�kQ���B�禸L}l;�zE"�a�M�H6~V=^3�q:���0�RX�a�ոfp��M��v(�1A%�<�G��GP��yf
da�a0��2eL��P�l�a0�j\b+�6T���;�r�#�r�zݹ�:3��'����;���M�ߨ00�%#���WazgC�wR�r۝�1�.a��ؤVč;kч�!/,�	Iv����/�0�Π��Hg����1��x��C�����I��6k�)����*Ge=|��e�Q�`ӽe?�gJ�&�mm1�*{d�VL����E-/^Z��K.�-�V��d���%��[�SB_w��S�)�J̠�="<W]��ع<�+{|�b%`�Ii�ׂ-z�"�,���5����q[�GB��s���
��z��q$ ��#>��l�V�%�(Z�س���S"�h�ըH�^���[|ّ�H٪$Ђ@�Ơ�/��}�tp�Q$�1��U��'_�3�n���basϬ���:d������x��QnO��^JM۟����c�ް̄d�M��ٍ9����A����e�h�F��}���yM����db�3=��������C�e11��.����d�n�58�y��f�%R����]�#�U�ٷ'^X��t;��4XW��t ��t�j�4'����YD�O�.���h���Tdp&��|AY.��ު#.{�E���p8(;����XX$I(�s��6T��nfB&��w#.`	���3��\S����*L���$��P*�}ׁ�j�Yz0��W�đMPJ<���7�^�=1�(�(�x��Zՙ��ڷh�˴NP�s3�Wj�5�1��d���ƾI��w����� ���6��I]�ĳÜ��)G���ِ���~�HJ6;�:=�2�Y��Թ�ߌ���O�ܸ�+G�h�R��� s��M��؅�� ��i��S����7�v�d����Ç?)ғi'�?s����1=ś}$���g�>H<&�'/�+�w��d���ٰ�㡴�z ��A�
��V`{��*��h��v���\p�
��,w+��9}��h��+�ia���cq�H�4:��]��f1Z��i�%�`�|��Ɛ/��ۑ#� �8]�_l���9D��Z�oO�x챍H����H�AE]/���kz�ѝ6k@��/u_ς��������W(xPBc{m�6����V���U�,�sR7^��r<ɲl4~�X���lů��#��f�1�ř����֧���g��m��(�4�f;�+5�%�;	0
j�0_n��pyaF`���5m����W�L��xmKLJ� .��@�H[/Q*�)=���^TeZ���6l �<Yw��bOh�֡K��z�0(
�����[H%mM���5���$���&Ʈ�6�9�A�����t���" �H�������$y��9�*�+9��%�ϓ��)=���D0Q��(H��<��䏄\��������@T��m(f�56_�g���YR�P���L��]�_��;������c�� (�7ЗGM3���J��`B�_Y�n31�GI��βY���eCM�ٛ�T+��$���s��֚�X��[�Ck�`v��'�&2��	I�9�'~V������<��Vˠ��@��/e7B�TW���.&O&�;�w�d��?�x�)[~��.��`��C>4�7��c������:������O$_�/������񩫂s��GZ���wO�p�o����~� ���2d���-�3cli���Xk��D���d&ʪ>�[��5c`#��5u�)A���0���6g1"ͲI������M�m�i]�mw]�G�[���X�7��z1��!G|���G"��-��1tK��EE������&��Ϋ��pn��p��l@fV��uwm����)N����V�@�8,I8�������S��M�=�C�'�����|Z��ԇ����L��K��an�Mo����)�����1������+&�m�pf�+���+��	���X"�c�}�h	�R����	r �z��B�������[m@|´7 ��\wWIߑ������ظ U���>xS�3f�	�ʏ]��<�v9�����| N%�7�/�u��)�$[�M��\R�ގ��"���w��&*?��5n������f���T>��z}fy�-��L��ِ��K�I�I���f��<�9,�]�c�w������iH<���s�[w��w�qp��@�,<g�?_P�Ep�zN��q�C�2j��Q�܌�S]���z�Dp�Hf�gk�M�Bt�oa��7��S�g���sm�S��I`����l�7Z����뾅���WJ��ҕ���ä)�!g�����[˽l:����#D45R"���Z�%m�Q@�o�}l��P8�t���@�ꢻb?D���������۹ߑt��t�^
�2���a{�m���I�ýw�<�j�(�L��S�;�@���~��:.��u������ە��i:R�qL�!�2���f&���_.�����٪s(o��\ }tm�P�-���l���f;9��������ʭ�tû����ݺ�l��������8Q�u��L��u-�k	;�����3��A
�R<!��W��ry���z&f���|������n�L�B��l�t�Nc�q��_ෞĬ���O�T�D.�隘c�.����:�<O0�0�C��;C%�~��錯�����iQ`�mR��V*x�B{���t��2Tg��y:]�|<�)A�!P�1P��S�O�Mp�o=0��ȉ'$cX� �:�����}�ˬ�(q�vz����$��������|��L�BOo�	�0H��~G��>�Qyl/�8���A`Æ�k�t�|�<)�^N�<P)I�`����c��R+��Tt5����u�� <J	��
D�Z]�x�3&�9?F�K�f��q�����Q�V��� �4"H��IM�W���\=L�-c��B�9D���M�xv!���D(�f���!:�8���ES�v�q��ɦF3�o���6E�ôe��oh����ݿ�Mo�+&G�.���Ð�����:�}���x�~��&�6)_m�lvZ$���~GկJH7@_H�SؼoW��zh�f7���5�sL���HX9*�[��~a���a���Ѵ�O�
K��gZ������CS���FI{�p�_zG�h�PmpJ�H��dU�7�o��X���f���u�/6�6q�������f�i]���r�4�\�U%@�G.P ���0"Mtw&^��\��-e��Kl
�k�����BV�*��f�v�N��rb�q��R�M��ĥI���h�]�_����zw.�v�>��O���p���A��(� �9v���n��g��ϛO\�ο��oo�:�w{�3҅�'�9�j�hb������\��~g���f�?��M2��Fc�B��������@O���J��r�s�XT����͗��M�'zN�Ե�S@�zd*�1
~[v��j�x�u�i<���ߕ���|�Z�!ð�i�bϗ(cÀD�v��H|{�����mP�#�Wݙ���iq�3>�!9rl��2�e�,!B	�޻J^�o6�_ ���g"�Q�s��	T������uь�#�7����*�V��%��1hPce]�m/j�a�*�����ֳ�t�F����c~�e�!6o99w	�$�6�Y����eqw�F�r-X׳T��J�Ğ\�pXF��m颎J[9�"�LФ_g&l�`L��c�j��F�^+�*$�A�7�)*A�$�P�D�x�r�"VX��(L��JK����R����)a�`=X�{z��н��kA�7����W��9H�R������(�:[�f#�ZG?�"�M�r�]-��IQ��V(�!c�<�ks���i��j/�'��蜒�L�������{�0)c� ���2����!Y\�(22��ڔ&Жw2ʧȭ�5cϮ\���Su̎��}@��5�"����an#@�"�l�^9X9&�1UV�`�P�b[Ǹ�t�\���~x��Au�@j�G����yt*�w@�W��ۄ��q��j�E^��nN�2h�� Q�p�,�������<C�oJi�P�E�	~�H��w �ʹ�U'ο���(���:��O(�d��rP��l�jt��z��8%7["1��@�ZN+�J�����ˊy�q-�k�>H_ �v�>�,7C��2л^�n���4֔���T���2��_kI-G�,��k��WG�Dǜ�N��Q�%��,�Z���h��RY�$*���1yy�P͚������e�ܿ&B�h��N_�"7A2�f/�qxL����Kz�?�VKZ�M�����e��
��S�8�[��M�4 7��I�:�2Ĕ �NY!��ak6�
��`;4D	���S�2]�o	�Ƙ5�:F�[��kE0+{�j%����v�ը�3��?z"%�i>7g�B`ɼ�@�g-�	j�D	�����s�2�l��$)%X ���E^fI�/�V'��/�O�۾��9p�	Nz9���v����j�|	����{v��>�Ƀ%PC����\R����~��6�����*��d�!z����e����7I=��J\��l��S�B�˰�+����cf��"��⬈��l��r͝���?�Quc�O�NԆ�o&mPÄQ#��K�|�n0�#ԩ�/M@�Mg�;����,-p�׻�YV��=@�#���c�D�G��!�kt�*���:����H����ª���T����~��["1i�WA�Z�� �+�a���O뭉�<0lv�MjpHf�s���s������\�G��<9���bߓ�vY ���/Rn�s�V
P|��/j\�4A���a�G�.q��%GC-�'d[D��K��4���]�d�b��:_�A.�� �@�x?���S�g���y8����JL�?6E>L�ĝt�飴��'�.�����hd��6�O�]X1��WE�qɟ��4D<l��v�ݓ�D�`��	��}zd8��`a[]��_j��ƮvF�_z|��v�iU�X�D�T�ݕ<1ĪQ�Z��-	�F�:P���$�;d��.�0�J���O�(4��Ul�~���3��	��3�}5���a$��ot\�8*I�}F��=Bkd\�����~�w��v9'O޼��E+�WM�����2����������V���y����� W�1�s.����Ϡr]�4@���\{�1��ޤ���|�\S������coiH/%aF�H�u�A��@'���`w���h�z�ؖ���������o%�Î(�Ƿ��H�6��9��\�j���)@�-���7������A��MJ�"mʷ�]0�q�O�����W�Z�&qki��!�q��u�8�Ip�u��@'lF�B��f���܎r�U%��J-+�H�L������5�����o鑆«���r��t��%QDF)&�bt;8��B1����j���M�D�f���*Du����ڦ��љ;�0�&JM���*�,�Hĭ���A���[�zI�$��|�R��އ�۴���Bv�T���m;v=N� ���AV]�6;�ޅ���!<K
��}׶^�Ԟt��slc�*Og��R��B'�Ħ�v7�J�F��{�)?�S	�	�r�UPr_�Hh�j�5�l�B��)�v-x�����Xo;����7�����ñ�~˘�`c&ӭ	�t3�р>��ܷ�,��ґcӱV$�t+3�)<"���'ӹ铠�^�W�+ތ����8;��b<��������&����G�t{ �M�ɝ�}zΧ��S^��p���h5j|�[�L�5[��]����б��m� �%/��v�_<(�y"/E*���d���k�*���A�c�^����5���Зb�����%:z@G����y2Xk݈ZL�GĒ�"����O$�4�-�Q��g�Pj By���%m@!b�k�����@:��7�7?*��v/$�Y5W?�j0�AO&'�Jm�\)��L_[+"sjPo���m�:��Ɓ&����	�;��uw���wJ��\��]��,�\��B����v��ٯ�b������T����8d�Q��2�˪L���y7f���TeQ+�3����\I7����ڭ�������vxǑ�Ć���f�;��Cjv%�A�B Bf�%��M�+{�9ᐻj�����߾��'�atb���u2,�j�"X��@�m���a}	-~�EC1	"�g6��
ҟ�3��M8�y���)�+<'+[�ͭe���+g��$���|Wpp����لE����Rb�B2������W�"�����Y#�W�%���~9$��^��t?��._K�1}j�y��Z�t��%1"� �^����D1�é��2��۳�֩T���잀�03�_�[S���>�%�:�j���,@L��r/�9���r�P�.E��m��X�s>���r�)��1ӆ%�!Z$�	��ca:�[���
ֳm��U	����5�d�§f�WYu�݆�i+�F��A�Nc6?�H�5���)s����Q�yE9�=�s����jH��)*A��w�%���v�+���h�E���ls`-sc��� 3Nn�3�/6@�jϖ)��M�qT~�dJ5T�FC�|����0�i-7�M����F?���|Zd�����B�'��v�a�<ø-�+�5t����Εi��d��q�����g����Lz���}�[��A6Z2�5��R�_�]����	y#���@oTv�<bR�=�ܚ��7?I�t�*�S]�K�%
3S��Y��u�6�o�:�U /����-=�1��F ����g��_�lQ-��F�XucX�P�` N e��״�ҋ��T	t~ң�?�-g�szay�.iJ�3���:��u*���C����N�u�kJ��)�0Xܠ��ԣ��%(���ӷ���	�,뺱�ඦ�K&W]�c����F/�iق�g�h��)���q�ɖ�9��M���Q�����Rza,�:�5�$c����w�k���@�
����3�u),r�Q�q����T�=\�	����K���=�@�;����sr��N�����d�/�G$�Z�!=���Rz[k�?0����%fP�l�է2�D��\�M�$�YQ�\=Z�G}��� �z6T��+i\�@���v��7�p��!=Q~�?�T�B�@GT��u�a/��BB�[�p[P�F��k�Q�T��;#�����#�vI6�����25��"�]��&���"�����e����b�7�u�Mw�=�-3�ȵ�56��S�^bU��ͨ���Ɓ�4K�r��Y��� ��٧M};��;��|nI����1��b��e�����pZE�K�t�-C����RT��|��]5pl�r��ɺ��J�:�9��Uj}������"5L��V(�6ށ9��:�i��Z@Do�眝�k�p��
�lΰ�)�0���(�0� 7��p�Tb>�)�����T��B�-�� �1�xUO��M�.H0�,"ĕiX¯f��D�ji�~bݰj!�_�3`*��L���iL;�Wz���cW�T�~l��C �\_%N��iZG���a+�:��@�wfi8���^�2�B��a�r ǘ6�US�v/"���6H������p;䳤��%t�%�wȬXn�k���rY�o�e�����M���j��;$�%J�Zu���d=�(�J!PJnm����ҽW�r�%E�����H��Ԟ,�}������+x�x���yQ0;	h8e��fW�������Բɠ�̸�̔3E
hkvθ�97zE�7R^	�-�#�z�R���KZ�k����}}(�����*����>�tWm��`>�K��Kl��@I�⪅��^J���Cj�V)��/���-�����e)�������u�)��NZT��pF�l�(�=��J��$�����2U�~ՌĎ��ҥݰ�d˚�L�lt�((M�Ӏ^]�P'�z<�gdX�Qg�8ax�!S/|���2c`��-d��:��>�q^�
:��s��'��r��n8.�ˌX��Ӕ�:�M%����ȶ�Sex������81���%m��g�ܥ�Ob����p+�U?+�3�Ƞ��`��7�,{^�Jf����8����a�5zY�@/Z��t-E�qQ_��d��%����
����ڭcv����]>7"Ź���P�4<���v�R�2
�i�X�L4��4�Rqj��򯲖�0`𗘹���~�K�jJ��f34�P�ҳ"��#ij&�z/� t��,M�y:�Y7�&�^�Lt��O���G�u77BQ-�Ċ�F�3x8���s8�Azt�����������ʣ��&;��e����<WZ��h���}�&iA�z���$V�9����3j��rg�vz��OF-{ГA�Y]^�F�Z"��S.�##�����7>� -��.BM��1��/�?p
����~�O��m�B?T�)8��Ͱq#�Ȳ�-vt�l>������'�ު���X�:pm�?�������+!��T�T'��*L� ���>Bg�h�@�܆W�0
���֙n�;�R5�w��y3�Py�����@؂%����!�&+U�D�	u#��K��>S����W����4�e�N:W��R}g[x?-Wq����Z��0�}����L'.�WcS��"�g�"S�+�K�"|�⌳c�����,_ڳ�j��Rq�܎�ϩ����g�T�˹�Vi�'�#��?`��7a�#��#�Q��d��������#֡�v4󬈲����2>C�t">o�=�W�9L���L�s~P8�����9[ &O�x!.�kIBf6����R1aOBL�v��/��GG%_�:2�������竏�g�(���T�,H�w�C�!�j�tO1���oLj���Mk����)e�e	m2��n������۴��£�x/�1#�B�5Tt(_�eT��7���4ѿ +��!jgP����N�&,���=?3kL7[|��p��rhh)�.!Kym���{��\��ۀ��(�V��Bz��B�A�
��;�~���b��}u�5 �[v���o����IYKW�����w��*V[<ɡd��-��~7��M|`���D朒����U{G�}�x"��r#ܔE}돟h����$�NB���hu�������y�X�{��oW(�%S01|}�T0i}��N�G����� �r�X
�p5��M��E�<[���ǁ�?6Xd|;�C���K��trsȒ��B�m5���I*_
�n������` �Ȇ`��i��A�Hj����3;��	!Y�۪����\�኉�I�������� D��Pm��Bbo�n����p؂	O�u��k�q�ug
��w|�0D��K�:�=����%���g`M�:���W�S^�2�
̤Y_mb�8��vѲ�S)�ZS�;"X�R���b@�F`ٯǀ�����`��3�-�\�9������4�s�N?@c��޽�G�Q�Vr�M-h�y7�_��юIQP�q�|
3=�K��~ �w�]��:�:�iD�9�	5� QCm���o2е_;Ӫ��K��23�|���Q��(U߱��.u�"��_.�%��֊-��k��;�f�c�2�zŝ�����Pb]����s�������������EJrmNܴ���<��ܔ�F ���r�T���M�����ޥ~Al��%����kd<j��z��N�������U�Y�L���d!3Y[M��	C�UW�[�eF�-�(̅���E�+`�r�<�(s�1-���U�u�t�AI�K����<PN��S*[.�M������jQ+�������}�e�dhr��LC7