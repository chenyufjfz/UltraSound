��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e�	X�Dy1V.Tٵ���E�n��i]5�h������5�xA�� �d p���h�t�?|�q����b2į| ��ע���8��:���y�HO_����T�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬��q��lv���~6��kU����S4v�ѼO�4��\О�S+�]�����2��@ﻤ�|h�(��|�5ז5�n�
�(V��E��pwlj��p�	*)G���B�������!�A�qE|�u���+5:���I�/���ׂ;��-�jP[�F��T+�kt�/^ϵ��2~�:Ǯ�Y�F*�ȵ��_7�=Y�"Y�z"
mWyɞ[p��q�E[�vj�L��В��W� nU�N���ӭ
�F�{ݒ{zW�#��#�Q!�7���3O��wV�~�����F-լA�w�/�f:e��eZ0�i�d�ư���n�΁z:kv����x��[��8�ڂoI��]�6$�a[K�l�{C��#67��l`O���g+��6��m,��?/���0Yww�Z�e~�/Un�Om�&^y��ց��b�2'��d�����w�������S����-?�,C^iY��10��g����,��WhоKt�n�ِ�+���/����
lS�k�3U*O�<��ޫX�Yz�-4��B��R�33�Y��G*E%��
�,-Ԗg'�B���>Ş��Y �?�}S�@b�q-��mBth+�f���*��Q�B�Ρݼcz-n;�ʵ��s&�������$4�K�����+I:���4n͞�Z�t)?X�8m����'�J,�?���LD�q��>����c�rC���wj4 �^��0�a��2$&�H�Z!`���<noɖ��Y���-_��¸���w�:=�~a�|x�! ���O ����!����Bξ ��ᔇA_UÉ�7�Cp*�:[��D,��� K���K;2���G�����9���`c`� 7���L��9;���"����?�F$�+ih��ND�9����2S�r�??�>)�)>��Xma������iǧ	?�@��H���8bު����R=�]mI�L��e�ܳ>��o�zjRjB(�F���T��+��g��Ɂ,��G��:�QJJ��A����
�c���:M���F�>��Ir��HgdFyk����kI�Y��%�k�1Qw4x��erVʓc�e$�`��h!3>E3���e���o�)��g�2(����H���mYE9�'S�y�&!&z���p[�MT��#y�Q����a���_�O�d�Rm�2�)����Iج�}m�� ����D���0/E��d��m*P�	zU�X5�99/ʊ����"k��*Ak���p�cȱ�`N�g�xo��lO����(�N��	���Q�j��ڇ{�+�����Q�Pp�7�:"������>?`��#!�}?u@dQ��.ޥ�֣��1'����.8/=��Q��br��+xR��� �"Y4/�_/k3�e���b<��U`o{����,� m?�I�tDN��$�8�:S(��k~�* /�u Blz���n$D*��4�V4Fzi�q/���$���zEl�,�ف�
�Y �G���;'�F0������\M4��N�f���^
t�?�#��E|$��m>�[h�1��$�t'�K�t�{�md#0�z�^��~�w��F�o�kq��Z:ik�k����%�!W~g;Eu 2�%b����)�^�ㆳ#��#�ʱ�dq�Ú�*���*{�[�Ec^�D<�5�_�-��2�Ƣ���Cr��/��Wo�4�t��5�����=�s�d5��OSN_�]'J_`��%��aw������~ń
�4>����`���}fH�YQ��m~��Ņ��&�h3�=E`�)%����O�@-[%�&��j_8����>����{�:֩4��{�{������Is)�#r�a��͌��{]8턛:�%F�.2k�`2��#j�Xe�S/!��ט�3��k�E 4y��Qn��(FOY�CÛq��b��5�a �K��z\�6�3�������Y}����t7)^Zk����#T��K}O-a��;�EV�*W/��O��	�������X7�	�c���[gs:R:9���>V�ш��nY���ە~<�<0��R��!Y��dīO7ૄd޳dU�W"�{)`�]M��A�0+��2�O��� B|�QaG�P?BS�u�Eu��?�"�
���:��I�
�#%�Do:qŞ��3~�����,��d��X������w����,�ذ'�T1ֵ�i2I��&ebQ~Tև& @n8�m_��fc�I��}����D����9��<lg��#�*���H�,~x����o���B/̺X/3��l)�D�o�]��#���L�C�t�[�f@�,j��� L,?8,����^��X�6�'����z�z���a�v����/�d����I�j�2��:�Kb�q)���Sb��&��=e7�+�s��,�ʇ��ޞx\�ν@�꼦[�-���A-�|	��fi�*w����
�WuC7j�_� ��r��Ao�?�G��\	�;��Fg!ɗ����5批k��]D��z*>UY��t;�<ڨ��P���[��u��Ҋ�q.�J������\>N����0���/Y����ݞD��uP�~����s���w$��<v�GT܇؞�ee$�XgkrW�-��)~���:��i;��6Zr��S76g-HcRR��l��X�������t��s�m,��gR��7X�`�_��Y=$��<q�Ƚ��Bz-��1�sz�n�=5�#��Ϙ[2L�7E�>�,w۫|���
�F�B[ ( y�3�}��P�¡�P
B�-�S{ȬY)+*�(�' �Gл)yGp��t�pn�_uq�C�� �	Cˈ�t��㗘3_����vI
�#�~Z_Р`��Hh����~&]bC�	,~6�-,�ePO����<��X�l�B=��p�Y��ֻ
��"=Ľ��u¹n��/i��]}�\峣�}ˮ�j�
@3]l�u�@�s�t���&D����գ��:����iy]yZ�$�-(@������ZU�*�+0
u��HI���&�����sH�>�E�(����"��g�M�J(z����f�J:��Ϭ0�Г%�.=k�L���6�ApQ� �*�#�}�u��������=OC�e�PO&8��	��覬Ҁ�d�\�������P�g�:�,7oPp�׻J�-����=�c���-8����r;�E�Z�<|�� C�@�;�/�lڦYd�e������i&���<��T�}��f�3�>�=E%>�8�c��[��F �N�:(��ȗ�����Z����cۦ��t�?�R�[�#|��r�@�-9��9u"-���e�����MP��A���R1��f%���.����I�˰���t 7s'��e�H�DW&��ʝ����;��<Vh��J���i���Fy?9�y!�{�I�%%�Y��^��3?vM�.�C��a�!��H���ׯ�D]�y����ZO��n6���QC��nkdgjFY*#�#�����p_J[�"�_��:)b�SM\W�~��K9�E<����{�����G=*���wk]( ��-��pC;�M��w�҅�[����6�E��:eظ�e�H�f��2�ʽ�����ː� -�:��P� C#J�� Z�6��v���1�0�$/��N$p���f�_UH�u�)PtI7�6��RHG���O�B��%�|8��Ov��STi� ���>�)�����~ji$�`,��G�b�M(#J�=`���=X�z�j֙�K8N*7�?�_��0,��W��#�02�׺��4o�-�(�<��}	Yh`I�L�����~?���2wǤB�$�ɣ�lBz�C
$���	NI9u�ظ�*V>�@<���7Q�~��:S*Ǵ��L����랪�Fb�ᮼb��S�p�&ay[VH�2��i�U�&��=]�3\9����q�%]��:���%{��<�Bش6��=Q[tZ��q�f��U"���,�a܍�y.�{�aP���(��>ȚK�ZϾF�j��nY-8x�4���_��/���`�����W��O#RТ���c���<�/ys����[t��xݑ���L����P�]�V�`kL�B�����\Ꮮ?��0M���6����M+�h"�ρi���]����S w�H����F�ĝ�
�c驇��OZ�2g�G�;��>��#�U�� �:~F�J�ioT]s<��/@2`�?�t�R�]lT�˅�4?ϙ�7Z�֎���#�Mؗ����^%P���W%|�Z��	��^�(	#���AI'�P�)�D����u��H���-`�۠'Jc��QQy�sĺ Հ#����>8>'ʰ]4ցI��?�	�	!;m������yw�Tמ`��J<^�^# 6Ǭ��5�k,WL��\�$p�߇�B�`�4��0��5���J56��$aeC��������s�"���y�%�qE�v/f���<ˁ��!H��Co.�z���N�,$���D:��ص�0�d4����Kf�J�5��&"��9�;F��1�&nY���3�o���{013c-��M��Py�J�K���j�{��MwK�ad�i���"�!m�����:�������^̫��
�w��Ts7�D1��f�՛`|$�dUO����vt��ER4����ZB1I6�e��7���m��r����Q�� a��_sU_JCޒc+�*��@IL�/&ճ���Fh���+���f�F��a���o�����HE��)W%��K�W0����C�_ӂ��Z�N}��M����!����:�_;��Rb������l��Y�åuZEc�~J�t
ɝ} L!�'�=9�k��{f#t�p{fNE�7re0u���rӪѺ&�U�m�4�.��Coa�Cz#Gl���p�5�W�[���T��xi�,�Ru�1�|�U�s���؞�p�*�|*�Yӎ|���:b���R'��^'��QG�ǳ3' �᪉�r]<9L���t��P��7�� �3�1�����������y�w��Ĥ��e�Z$���{b��6�,�6a�ۨb��t=������b��l��.��F�O;�"y����P(�
<uj��>�d-��'f�d�9m��ҹ���|P������F�ػHl�`@��f�;~��ΙR���$H���;�[&֫Pc+���-rܔ��%�䮖�*k�ʷ4S���x�KW� ������>^N����"�<���Mu�&S�6t�������V,d�k"r�Q쯥�^�����[�Ͳ{���|�oCN�CB�ZpM>�:�·#F�eP�� �n9�t�7���xdn ���3ݙ�0����Z%1pT�DnO�����:�-���hB�ʸ�Ī��p��H��^w�+���~ݦ��V�w��� m��vG���)��r�FaVx������ohw�FF4[�����	(��y��ԟì���h�f�%�jot�mC{Va���A�;�:ik�_�U��%VF����e-
\���|��͒�P��v���pvE�ڰ������f��q�o
i��"o�;R���M zG;��<�A�޶��P�e_�Dۼu��5�/up Y+�yȴ1���,�p�.걉$0���~�֛#��0j�,Z�:\L���J\/�g�@,��b@)q���V�+�]�a��J3�f6oܑ�	�x��&v�A�O��)��"�i�+f��$<��n���{�v:��h0��'��އy�����p���y����F�o�ѧ���v8k�z���-�=�����őe����IE���Է����x��0e�h�YuD�����ڮӋ����ݩk�tl��F��sRd6�_�,E��9�"s*N�����M�2[Jl�����	��b��Yq���`|;�	9�9�Я�Z�6e�U��4� ���!�y뾔���ڡݝ�Le)I^�c\4A1�����,�s���f�\X��`1�o_DI��0�H�.<��ڻ�����̡kM��ZÜ�lX�[�����4�e��#"��<@&��6�?�ՒUo�"#����x\�~�W��A_����
��a�E0-_\Đ�M?�4�(�j<eZ���'`�;�'��%���+��gy� "�*��8��>X��-�y%������/�d'Sk/�� �E��&��i�kG�*}ۈ�u��vxON�!�f�v��f�?�c��dQ�l�������\j�/<T���.q21�YƩ�����.�uN���o�=8�!����GXF�'�?H��b��8�:����KLVv�<H[�O��/Q���OZ\t�j�|�[4J��hG;22�d X8�i�?�SfM��E�q�p�il2�ST�~R� ߱#tY�v��c��Z%Վ��S�MT,�$�����%f:���:�b���,��G� X�=����s�������@�.%(���L�V����p�����ek�n'�<43�[em�x�	�UvOF�'%�(�7
����e8�&<[��A6T�z n�C���@��G�
z&I����_vO�F�A����8��F8�m��&��o#�����ӽ�N<�	�'�н���PpK[��"#m��:F\�͔��$��]"#�{���:�{q"&�jY�l��U8�=#�>Ԛ��l�����$��B(_ɕw_��ۓ�&�v��Q�*��f��p���G>�B���F-��P����=��+�;�_
��>x�5׸>7G
�"�1�,?��%��?�J�u*�.�@!@Mn�V���� P�������e�c�ڞV���+�-˫���Xk��|��}P,Px���>ǀ�%ţr(���T�\O B�=��1[0Tk��d#Q���-́)���1@�B�1�� 54V[R���O���2���Bъ��fM�A��ŋ�63�b�E2����w8�{-����֗9@}q}m��J�G���'�-y���^��n�v�xF�liP���G[
�4�\�"b��=��$0��s&o��KC��夵�k���#�%W�j�o�/��ñ1�V*,�4���m?�u��[���O:�;6���PR*<��!i���)S���W�e��� �7�䃚TL�'I�V�a��^&\eo���J0�����������Qł+��0¨�Ǟ�}ed�I��=M�w��	�{>���]���c�z�e��>RS�����k/$�_U��̯ޓ~mk*,�e!�/�����Rb={�IH:Y��<l(�A�Ȑ��eؚ\��Z�H�81ԇ���^]W��F!Q���4�i�~��]�Йs��o����b2�Q���0��ʛ�{�%A�/&�u�}�}<��=�	V8�{=[[�aho��)JS	!�fD����V3<+˂��M?��;��뱯G��봍��!j�bđ�\��E$�A3oF��#��
|JSOU{+6eA4mÈ�+�S�&�d��}��.�CڕĂa��״�B�2dc������:��! U�^!�0t!�2ҷ�,)G���%�7���x�y��8\��QS�bB=J�WN�p6��"^�e�4qr�Y�
�C�e�UV?g{�i��S�L��i]Ŕ�ٍ0�nkn���p�<$~��hK��5�8�2�":~L�<�Y���s�R,�4�=`�N��Q�I8� �Y����MHiĳ#XMƃ�s�[=��n���κ�6�$�Kq���VQ��\o��Ҏ�i��AӋ�~�W�a�w� ��!5Mܫ,�f%}�c<�;6�ս���;4��ȫ_�X�>(,�`��D��ۊ���;�D}R�	��?Q�?OBbH�V��$�r�o�)��v#�	_o�������QK�Y��x2u��M��K2c�v��e "}�cL㉾���'u�~����P��I\�8V do� ����C�6�;����2���P���G�һ��B�D���䐖:��Ϳ�xt�ϙ�a��ۈ��ef�Q[��F��y����z�h(�mC�1TX͙���j�ו|(����p��e��)^���)D,�+�ڑ�́�W����˓�k�X�|� g,�` ��`��3]�/65;%'Q�2���[�׸|un���PR�8�(�#'��P�<E�f�/s8i{�N#IQ���X��QU|F���Ks��>u��������e�"l�jR�D��j�x���Z��nM�`H�Ө�;�R �0/��i�:Ѡ��ň�r�2�3�|G]_�u0΃#Ձ��ʥ'���wjw(p�]e�2t}��}fO��o�G�
[�dcL~	3����-.k�/"%���q��P���|��Ѩ�N�u`{�h&T_�^��]' ��y�5Nkٱ�K��'^z��{
;��H��#�,�7(<�����D���w�[�WG��y'�{w!{;u��@��T�	�ʢ1n�5O�~��׍f�/	P��o$���iI�~�S�C}�Vz�o0�q�_��A(Z���5�TŢ����#�ݏ����}Ԑ
�Qq�τ��v�d�Ӯ���=͜�Qɝ@���3ݦny6�7&�4�*��G0act�3��ci)=&�e��J�2�"��(�T���"�?$���{�E|5�/�$Ԫ��1�f!�����o�#Ì9���G������+�t�m��E�+��;���-Z�Z���*S�e��)-�,��z� nc^A~c�0A��,A^�+��TvL�e���h�D����P��6��+yާ!�+��w��j�p��C������`��P�Ez��&�+N��'��Z���R��	V'\F0������Vَ:Y5��'5m������b:�)�)pwW�ܢ����G7v��pȟ��-�4T��ڜ�}�bC��'�� �Ϻ�q�5�Ս�V_!��>�N]�i�Lo��a��fGʱ��!��:�Q�H�����F�v���g/�$N��'%V���||����Uwk�������ˁIK���Hxoi�MyM�2�������Z�q~9<���|KkP\_���]�py���}\�����i���	�i*+��w	�{���z������Kz��8"�u^���HDU���D�ܥf`!uZ��c=ӟe�`e��r�3�ٚ���4�m2���V�qG)�WRW�+O����nF�����=@ O��XZq)��R�8��p�7��(��6F%y��wlbF|ܻ��+-ce���
C�>������ �-��	�V8r]�V��P��|ok�%����١z_���vV�čM	��-�ͯǦRY{��#��1ݳ������%j�Hq�B�y��F���og�w�c! �'|J�+������
�cl�5}�y�C��|w���z2�O�UV���)n*k��z�}V������0��¦5]>=�`�v�G纒oR�pG���5��� '��g�/V���-Ib��a��fY���1)�{�Ӕ�D�kfI7�v��g��� �ip���-�c�Z�98\��cI���FAA��f\��}�TIg���3�?��~�=uL8л���k>D3%���]� �d�(���G��)H>4Uo��.�N�����?�?�u�OOܣ)M�|$Ex�m����0x�ɢY1!�HE�Pf��2�<�7(i�Y�GR*.��6sl��R�R9h��<.��ÒL<C�?|.
Ačm��2����]+�a{tc.u*A��/ɖ��{����	�*n0ɸ#�s;���@�
-�=.�a�s�U~�d�+�C�Ja����S��ow0�z���L?0q4���]1���H�3,���ń���)�'�UW9�ͮ=1.fD�y�]	�4�[&m5���3wDl?�t�v�иr��gt���RJޑC\�Bȏ�̅���ͻ~p��4�bn��n��D`��Ѡ��{|8'i�g�J�H�J�| 
�ۨ����Y5�`ZD@��;V�
�%��˒����3o6󼞒i��/l�h���i�r4���<,�GR�@�j�n`�l)v�.q�Bi�I���9��H_zbz�ʨ����e5њc�ݣսF�%�h��'2�l��s��~�ut-u�0��d[�����~�+6�!	��17��Ҟ���S{�!5�I��r��+�b��0?Rz~.5���Ԡ)\�Gk�t���:��.3�:���x��Bq�K���kx�_��m=�
2���t�4�"c D��#5+z�������I���d~���6����H���=C3�56�,9��
�����N�<��l.�G偹�/R;u�B�\i�!��V6�$o�q ��ݹ�C1��N�R`5M�䮋]�1���8c�'>s|����|Mv���<��r�FZ�a��+� ��o��_�⠌*t��� ,b6Cj�]d���;�Xn�;S���FY�%[��F\.G��R`��1=����-��Ѣ�`9�h�@����a�
���cIVᮑ���_9��B��#��!Ȣ��TM��"�W�IZq��a{|g�ѫ��K�����+�FI�Ab&X�?(���V}"�/�0��ѷ��v�����?�_��\%n��OjAN�M!��J�C&��D�#{		
dd�r���~F�*�Ъ�u��ʧYcA����MD@dB؂	w�X���.����
E����*�j�P�=x|g.���1���ё�S�]��_��?s�)H��`�o�$��|���2�O(g�8g� .���~=�K��L�7>��l����֛�:�%�j���1N�
��*O@�b&��2�����R�~������~�ln��f�`V��Q���շ��kE��|,�,�u�<02�̑��_)Z�T�@g�P?J1�J��٤Ξ9I�K0 ����.��Vg�����d�h��u�r��Ng��q�����x���3$J���P�x'��;�=>�����WhzFG�|+e����E\(˂DI���;ހ!s��>�/G�j ���4�D�����7�g�&%^�p
oa��ɣ���=������������G{hF77��M�5�D$[ߪ��R^�V�wfp@9
LK5&��f�Sf�q�MD ���#uh��W�c���e�W����e0cS�$�i�?��{E-
5^t���'DET]>��0�����8��݋cT1�3�~A�XSr��jPI;�0�'>����tq`�<�
��m{\8l�=�|��<Њ�E�
�uB�'�O}V04��ŏ�ͤ��#�G�?	2�f���bU�\+�od�%�T�Ԩ��0�l�!�8��n�i
ul\<\H�{�Ơ[n0]|�O~���1l<<��e'�Lk��hФ!�~_�Ԥq�
&����	�tD����c`s�"��Z�͕ g�����?�c����gܱuqQ0=sd�]��g��<�S��*~W�	I�,���C��V���U�Eh��R�n�U��N����ٝ����>�~���|LPo�2��6p�E���R��Zg~G>4�^y</�+g�6����Mᤫ�^.�3:*��?�a��B*�K���p�3��m�����˯�,�}�1ω;�����n��RD��Uw�}P	Q�/D��lq;�TsR�<ӓ�
p�yr�+�VVZ�*@/�b�<ɏ7.5�Ӑ�|����\�5{�X%�"/J��,���{Z.�������T{�,xt���έ�z���+�Ր|�F�)�Os�$�D�7W!�g�8~� o*�1	kco�� ���5݊����7(��3���p{�]�C��)�j��"��ï��~�����G~�xC��ds�wo�VV�3����X���	ɐ��I2G%h���Aa���1��Y��P�͑�I�X��I���{���D�nᓭ�2p�ޣt�ý׊�H�M�M�T��c��#W��z�Z�۰L.��b5o�}��La��OK�'�D��J���̊�*�Q���篲},_%�֤F�R�b����9�U-�(�w9� )�Y8��T���Z�Δ�\�z����g4�gAJGL�|��bR뫸-����u�ё	�k���s�ъ�����rb�L�c͔�&<=:�x����A[��0�Q����xp���<G���
s_��;�K�Ȼ<Zv��[��a/{�����ݧ}w�沂�4-%U��n4�E��V�i,M��f�����?�w[z`ɫ1�Kt҈��/hOΌ�.���e�>�����x��?���8����Q]�o�~X��׏�yV���	1�t[+<Z�Tj�x���U�^����=��W=�aF�6��B�2�A����g��
��
Wj�/���_P�%�G�"?��B��N3 ;�m�ωG��зD[�1qkxu*./۝i�*�$tb�Q~��@[�@�=�����}G$�,Dh�Q����6{R����b{ �/�@��8'>47OI|e�p�����	�FQSfz�F��KѬ�u�7�Ir	r%��[�	�:v��@%I�qROSI�@�6�^ ���2��U3]s�ZR"��ui��@�����Y���'�����b����ű����J����(@�O��Z����RӴEr��l���\��<�������پ�P����L<�a%^t�ü�~�&
�i�럾F��.Л)sF���\�W-���4~��wId�NZ�o�b���@��L&SiE[i[���6X�WwE�ߞ�O.�cڲ�jshF؍r�̍����>���9�,b^�l�k��U3u�l{@��"�M���0�IH�٤����\z2֥u�_阸q��>f��f�RH�r#�y����J�
��z����I�H-B��- !%���