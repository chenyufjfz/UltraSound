��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^7/\�ǘ������W��O[b�^��nJ������`Zu�i�[��Eu%F>�,��ry��� �]�U� D!� `{�RK�ф�9&��nZF���(s�w��x��ѯ#�V�D�D������]ӵg�d��j�\ �X���SBN�?�&��~�o=i���	��n�����«��>Y�7�]Y���ǾW�S�H�������'qs�+{m��-��7PE�=���D��3Y��po!呻�-�T�\"�����K6���OMŦ��G�$��_C�p��%) I6� +k���k$�ϫ�ס�κI�~'5*�/�'���Qǘ���6������|@��[R����.;e$N�VݩtV{-֎�E۸�7����T�2[�-�7qN~S/Ѵ{����=��=���ђ��;k����$ڦa��D�Z�,�����4D�+Wv�4-,>PhR��������P=���$�#O�� ����&��mTm5/���稰>di��[b�������.c@_p��x�`	���d�;�uP��e�J�1dgĐ0�_��+K������.b���w�o[��<�v5_�*�!�mA%�2�F�~	B���a�a.y�*�c���ܡ�m0Zs���8��k�h]6s^�Kk��;�� ���y�!{?�ﳡ���xk�8���k4<��owdo�w�����%�!��afc��f�H�oP�X���p@j�,y������T���*0�"��8�8��2E�ۆt^����oj����y<���/
�ym?V`E���eq�L��m�b���/��q=z��jO{���t�sG)�A�a�)3Aeu�u�pq~s�8�=�T,ך� ِ��Y��(4�?9�pouv����{�Kv�?�<��72禲����y�� ��ZI?[r5���"o���1d�h�<�R_��	s-���Я�����N�E\[z�hwW�*���3�qx��J@��*	��% ��7Ը�����KA�a��Ր�u���G�π6~Ng������_i��%���S�]dHw0�$|�XP�j�&$�"Qe����� +}5�!M
������?Ħ��t�q�Yx=�9վ}477Jި����"�����х����^���.mQ�?��R}��?#�����xv�Yťl��V�g��]_*��\�Wj7��m̔?�����{��k~��j0��޵ ���#N���ǒXLI�l��_��d�z����yٺ:��U��i���L;pvSo\R2!nE�=��,�SJS�JtR�>YɾE��*�����6+/8�+\))޸���:�������7T-��-�t�R(�p,G��
E����2�{�����ocJ9���=w��|��*�$)�As��4�f��+e�U�hG�\��thN�qb"8�ktrdժ���YnNx᪱�1\�r������%��c1±�h��X�R[�]�m��wy�!����������_�Mз��.����߂,.���;���e�)�>%:gϟ��Q���nz�GH~�(� .�˘�Q�ʙ�mg� aάH+\�cV�L˚_%��(�?e��=5����vgc���+��h-�cN���	8f��r��U��"����n���fZ�>�C����'��J���TxZF'I�4��YlkP���2�g��C�,6 g�6�|���O��X�ޗY4	�A�':��/���X'/�������VL!g������'���n�5ɛ>�w��g�b��'ף���TA��e6�P.O��%�U�ho����6�}kצ�Qo�w��;W��Lk�R�(�䛾k�u�l�����1\"	;��/m�e���Y�1���>D�����֒>p���X�	���vٓ� H�MdV�+���m��B�׸�;i�Dd<!��h
�l�aM�&�jD��F4�/�~�h����R�\(���[�H�#4�R�&t�5赧�ˮPf�H�.�G��ޘ(@�_ �����<~G	�H�Fe�V�`�}���� ����ϴ��x�ǯ���3�����;V$����պ8�>yï��Μc�� R�*�/1��
ӫo�mAe�o�j��P��
y�����7Bz&�w���z5�׮.$�3ۀ�f��<P� �/�ԩ�sm�u	�:�Da刢q��aO�0�s��t.�$"t[��`�EM�|�������[����U��)�n;ils镙�1�)�VtWd�-ٝ�k��QC�6��_��6jg��W�䠆&����ܼk���>Q[VW��*���0a۪�Ha��38i�$��HƵ��k����l6��5(���#���Zq�4��@��r+~$&�
]6��,�v�GN O[m�l�{fsw�Ax��)���H���G}�O |�.B)�b�@���$�хҭGƠ!W92�k�ތ���\<�a00�Vd����+C��������/�V&UE�T�K���_��Py�*=O������e02L��p��؞�>X)���l����I�Oʯ=��ڣO�OED2j�*5�t�$�f�̪;n��3 E��a�;a(m�=ư�����
�k��*������3�P�%�����&��d:)U���s���|Jt�aL%D�P��@A�"�]�F�i��@����;�\����[��/������.s 1d:�G}�nK�b����kp�H4�?sN��K�e{ns�㴹!nwݩt`/�ܙl`�R�Y��;o|eN��
֯`K�M��#ZA'"Y�=����G�K;��K��Ԩ��,q�me*qCnub��l�U�H��#����1F�B*,��B�|��1�L[hDba��ir��!E��Y#n�1Xo��G�F�qY7>�f�(: q�����ʓ^O@��J�i,�y/S�y����uÌ_0�q��"ZHs��jXU��R�5���z�\�}w�ӵ���E��Y[)��o.�	��Akk��0�A~��[�5�f����;���IsX�~{��"��ܦ<T�D���QqC�/����s�� �DĒC�'+1!{�Pqw�7j��D'����n�>�r��,�0\\U밎u����;;���e��CqA|���?8�6����Q�ft���0��21�2�#��d�������umss��x^�w*��vjn��@�_�sN���$hMo��������T�Ծ2�3I`�S�=
2��Ec+	r�H��t�v�y�7ȋ7�Hy���f��9�*��z�-�B�����:8�`!�$��'�C�R�U�e�U�˲�]@�T�>@]�j�m�o�t��<F�/�;�ƨ�1�E�L��i�:�
E��<ϟ�;���&]:cq���I%��@���v�,��D��h�[��%X!iǷB���(t C��ֽ( My�4�� r�2�pz���I�ߝw�]�W��ID3���yC(�6F�r^.h�0�ġqD)��iG^��86"��a�A���p��t�<ӫN�::�%�I�2ٳI2(��#�*�k�f_�@vh�.�9��u��(	\���â�m|� �X��ar6 �(�`}oǟ����y��<�&�d��)��N��FH~7F���E�R�a-P��h��v_�1u���4�]���4Q��uQ������|8�/�>��4M�3�v� ��Ƶ�l�i�*{����&��)�s,"������
{��c������<Ѷ�6���͔6#1�+����ڥ)A����|��}�5d62�Qfzݯ��2Eip��^&��n�wm���.q���R5YTG�:.���O���d�tM|=�_@�_J6���a	.ݭmu\�� ����t?>���)��kgt��z�a�a�%�]���=e�i`Ib�]?�8�d(�ޚ���Vtȋ;��E�{��2�M���{�8`@�4�1>�s�@���&����UG�}�6j�5W�~M�01����<��~w�sy�EB�L�7�k�/�ؐ3�G��B^ݐ��)�8�d
�[�w�П�o���n7/B�i���A�8�&�*�y��
�����1�>~��XX���PCFΫ������Y�/o ������(���ArLw�ހ?]�h����%�"�3�-���-�X7۫�=�g�"���~�$�}V/�׸l􊀘J0�~��y�$|L(����zR�`��[�`��F|{GwFT	�yИ�?Q��)��jΌP)��A�Ew9�A�L�&������:�����o��25���K���ONCO��1U#r�s��Po�
ήv*V� �v�u���J�zhС'�Y�B�Ynp�ShJ�k!Y�f��窟��R�mV��h�T��m+��m�@�6Ӊ���7,�!��T.UT{��|��w-4�c)Ϩ[@�0X*N[�=���V�ŗ���ͻB^%I΁�L�C�3rP�1����:�
�]6c������������8����"<�=
ۦ	���wEϯq8�wǫ�'}����W,���Dm#�ެ���e/<Aq�<�DT�����r�Iǝ�<�;y�����u�B���<�U�x4�of42��; _v0<Ϥw��Pa��	����q4�遙_���s��v�H5��o���r�n�W����&��G��J���Иir�V��n�v����v�@_#`���Sϝ�ֹ$������o=�ӹ�ǯ�0��x��[��W��������Sl/�9x|_����ç�*oF�]BZ�r�S�B���{5�q�*�u*ih�:]������l��8�o�P������3�βv
n��J����g��IԐ�&�� �B��9=���T֛��\�2ds��5BB�U	A˺ѫ�X�.�
 �W# !�F4ĺ��U稑�a̻�y�#;�	��M��@��b�jrDC^{��J���Տ��Ұ΢@V.��3���CO���w�@a�2��xDq���DtO*8]�ސ=�P�����k7Ȃ���#\8#x�R�Kal�)�"��c
ˁ�}��X��\������X���c�)n[�'���"����N���q��s�G�$ZyU�T�f���<�V�\�I:�߫O�D���f�C])7*1y����N��e�ۜ�����3�/���|xk��DwȂ�����Y:�#�,�
��ǩhr�CN�����0|(��#<c���t7{Ii�zZ[p�^��jx�h	��J�����q�0@edM:�:���d�w��^:��H�ޛL���`!Vhd����	g����ӛ�Ț���d9�-�G<�2n��p��sV=� ����Q4f<ً�pڼ�y�EsP�jb�N��r.�����/�K�)��`���d@��]�S�s��>T�6t��,F�Y�n��V�e�/�QBus,*i*���r���x,��|�M\s�}]r���&�����p�^K���0�E<q�^$,���ƄD��I�0Q�oR+������p�d	.U>���_���,�E��Zk�_�)�y��ω�<���Kp���l��>�S��m������H�	�fC�)ϕ�c|�Lb!�j�+Ef���j�f]d"���#�=���_&a&E���,ő��^�:a-�]��:�}*�����P%ElN3��ڳ�����)c��W��+i1;��]ك/k�X8��A�Q$g?0,`�]W�wvÙ[����p�I8���PNu��3�}�-ek�cx6���3�C?9�� �����G�	��:� �M�D0x��Ϸ�n�~}B3�D�􆟉N 1@��!:��?���g|(y]�gVql���P�5K�RfN( �6��D���KN� �u���?��ݍ�s
Ť$�f���&�!*�g�[�x���P��؉�*/Ai�gK�ƮZ��np&P�A��`�A5&��=��̈��H�+`xc�$�&d�rhCP��IC����%e\)�fC����*ڍ:>mȶ;5p@@ou��u�e-�FS�J)h�O8hw���U4X�O9�^�j |�a����%�b(�-��xW�gXd��&�W ��ہ��֋��+����2����77J����ew���wt�7�� ?�ʤ�U�sv3��Yp������s�ؾm�Ҧ�N#����VW9�%�G�Nm֌����-,,�V��84��N�/�~�[CQ���-�W���Gp�؛�D��>i�'��Iw9�W�	�-'�ش}�<�x�kf�ޛ^��/�T[X�-�Z�z�p>P���X{�W��� �"�.<��sa� �u��{���W1�	��e�qaM��S6�7�q�Fm0�K���v����/��3�̐/A"|��܅/�پ�2M"��������G���5�w�|9��O���uo��̍�muѣ��B�	:����$�<_0�+Hktú��D(���*?E��>�׻~�����.6��1{{�`�\�1��0���Y�%����Y�q��,�O�p�/��R���pI2���#���/�|�ZW�A #���iy����o��E�p��E�L��/�߾{Q�ќcJe��4�\�=�2�u�%������tB����r#��&��^z��*7��
S����Ț+p��Uf;�ak@��%6�����#��K3,H����E��nDЍ[)�Բ��F�]�����j7�,�5��C��i^�m��v\r��G,|�]��Q����hY��Ž�7�)��e�+m�o��eZ)�����,��Y�: iߓ&��z�dK�;:4/�ؚ�R��T�r�E��SM3Fg��x��
W�����0;���<=bQ���S��8!7'u����<����"vx�<U�����1/� 'y��9����_��P�bsJt���$�2�V��xB���N���`�	��8�'�b^����V�4*�����ĒAg��L�dR�8ͽ��*W��`���:]5�#G�
�5���ߺ�"j1	�?� "����k�Ԙ�g�Y�Km�_ق3�jr�|��ٙ����>`[8\f��_Ӛ���@cSR��[�ӪW�Ŭ��aJ$[�UA���{D��ru+���^���'�;_a4"����491_�A,'�/t��
x��2(��.B�����R6�}{^�u���|@Z��@4ΓQ\�P�I��W[ ����)�R�Q����
J�(EX�-	�����b���n�V<j�֓�����ԉfoeN�7��əÝY[W{B��=��ֈQ��P����<�!oϜ}Q�v+c�3�L;��;�ll�^�\G��Ot�K�mݺ�^X�i��>Ώ9�#��{1�#���������"��a8KtI��)���N@y���Y��X��C�.�����<ģ�c�p Qt�?��
q���՛Û8"��ziߴ�tMGj�?)�G���-@3ˀ�i��F�� %�]��5�$��F��^W�W}��"=�������g������"���`���J�׉OL�M��I[L��4������;+�7gK����f�)��A��O6yɔ���e@kR���1A�N�m)#x��hʼ�
"��м�ܮA��y���8#��?����3�u�o��qe�lM��6��/��;���:�R�~~ޓ�.u��DK����g��&j�tu9S������"[��E��ζ�����u�4����$��Ů�r��� ��0��� ~��d"�$�Qӌ�J�I�:T�\"��#O��2����.tC�I�x��J$�JM�0)���L��7T`����|�E��㑅�gz�B�H�$�Vzӌ$�̸�8��7�N�:���KRt6�j���v�|c3�e
�O@�pƸ��+�PװM=�Xq�	@���u
蝱��^�|!�
����/f뽍��-��?bd#}���xKP���|�w���;R�	GN�ϛ>ZU���9@%ncX;T�h�G�����1����%2�A�t<
dq��&�޻GS�bI!��m��PK�HY�X���a/�`ą${�n�q<W�q�H>�>�k%�J�[Bw�$FĢ��+$x׻�W�/���S\~�c�����\�j�O. �h�S��'�xzM=��z�S8�=�*A������>��`sW7�	�����4�e�sP�0)?)�k�3E�$��35����w���E
b.X��'�����)�D�h:�N�<C�|�[QP��p��o�&@G ��=��E��\�������v�� 
�o6��j��n�?|�e�(&$U��;k��*τ|�-8҅;�����G�����׿�ba�"+�w�k����>��V� oc:GH)Gҙr�:6��C�}��H�I��N�2-3G��O�c\�N�r"0�բ�݉���rW��H�����B7�s�f��3d��S���� ��H�����+�_ Փ�h�������<��4L
�|��ޢh�V4�IB�_k?�!x����'c���\gu�6��O�$6�Uq������-��
\/������"���j9���y��bK&��[��o�����i��=Us��,Si#!�[i�\��J3���w!���zS�Y�E�2�)4�1[��
�[�����M2iqު"M5���3���s �D�2���\K�K3ii����ڹmCv���#�,�b��>5㼆0����,� ����P�"�MM���J�C}��圉�'~��g_��6�lg�؏�V7�_q��==�\9g�IÁS�k|�����h_&��j�쵁�o;hk)�cf:{L&(��`�D�q��I��L��a#r�,Ne<�7���r	��e���w$F1J��D���<Ǵ������f0R���n�R���O�bw,%ԆC���cqz��`�Y�p�;;Ӥ�PrN�j�CFB뻝�6�/�aV��`�<:(Xa�`���	Qcz���������U'6��{iZ[�`E��UGr$�����0!��m�X�>w�i��7�<��6��|�j�5�?�f����~�i����z�A�F��]���{��}G��d�����~�2tuc����+����u¾9uxwm�S�ďRҬ��A�������~�o�.��|HN[k�K}Wh�d��I7ss
��K�����M���fUI:h�>Q�2�����G�Nݗ�'L}����3aK��NۄS�؈o(���mn\N&��a1���T��'������+o�9~�A1���T�Hk)t~����\0���<"J<�d@��sW�����M�X���.�:�^$��_ü�����S"���`!j����*� �o0b�l��mX�����ԣf�yOlͺ��QQ+��,��R�f��O�����7�\�����uQ.%ѓx�Х� #� ې�)�9:�� �����x-6O�r�֋�ʤ��3S�t�~C�,����q?K�N�Ģ�w��!�#f�����-m��"�|�2��8g�ݩ�M1w^��W��ď�6�7�S�����6�,�S�����Z7B
|�i8�����p|�Ǟ	�-��M��5f.�SX�Z�̋�z,��@<�0ɯ$��~�"G�Ԏ/��Lbՙ
������\��1m���a��$��ϕ�]�-����0ӂ�J�=�*�GXW&�P�ʲ�rHi��2Bx��1�������X�y)˯H�g�π�(>F��Y�ś*G�@Al�kMj"D���b
�u�Ya����0 -7��\����I�j�)H��&����T���or������A*���;��+l#B�B���3z�Wt�̏L	լd.�.)!ܙ��Հ�j�6X�F�k��M��k�ܚ�8���`������f��ښ�1�wEXUß?�f~��Qm��k|,��& ̓���R��`L�#ߦȪ���nQ�zKtk>�$�X�+g��t�.Ds�v�C�����b?b݊�W9��	��2�rYq�{�X�.�.DS8�H�7�mU�g�����If�����ii�g�r�/q3v��E@���KC.�W���I�y���ۉ��l���=h�!���=ǇpQ�����A��|>����H1}ږ�xa\�Ƽ���Q9uX�t�G��h��a�y;�6tǥR�{���c�ȉ�G7˶PA]���v�
)�:r�,83;��<��v^f 5��r�T�=�)��CĻ��6FA�.�~#��{B��J��>	����_��ʽ)_�]�[J�|LW����Rd�����du�T�l��;�R��HAh����|�<JT��a��,
�
N�>���]�8��K{	��O�f�?S����g�1؍�<Q�XS!��`�\oOd����w��{�-s�8'#vf��ڌ���1����#�ëO�~�Q�8j����0�`��Xy@������c�j]6������VuJ�
`̀�L��\���*�
:mb�c_n2p��}�3��?jX��8�5nV��>h3XQ����hf���IH]�.o����e�Tx���XF�����B���8������&N��<ni+�$9|9��l}�yo�&y=�v�G�\sg3�ZA?��8��S�a�w���:��b��d�E!��6����`Єz.��]'O� p���<�X=����a{s%E�HI�-aY���<� tU$�ꌽIXGN1-�#{�!�Q:~;q��カå�� �p�h$7�w�����4�"Y|��
ǃY@ϚII�X�2<��B�㙖�e�v�����_���@4}��eģ��z���*])�����Э��RTqaYg�S�����t��x;��ɖ#t<�$da0>���{R�:� T%���1:cW3�������-^w�}��u,����Q�V[�����xa*F6�Bn��*����x��b8������� �Z0���/_��*#�2�*�`+���U	����*�8�˲{t1*�'Ҷ����0Z�~E$$4;-:��F6\�%��{��:qj��7�?�0�j$����k2(��O������7Y��?�z|[,��|B�RjW���~-�I�"�A��i�݈�G=����c'^�h�+-G�)Ln:����ﻹ ��fH��2�D-Y㾴��rM�*��vF�h�);U���|p'+U�7&��Q�M�~�eR��(��	�d����׉H��X�dn1qp��G�:��ѕ�.	�\�Y2W�R����x���k@�ǻ��PP��94uAS1Ws3�{G���p���RP�v�X��yG�D�3b���?b�i{�� W�Y��ioKe�g��j}\�����T��h�vEy�8H��j��QHǶF�Y8=����5}�60u�A�O߾��ZJ�'���"H:g���z��u^v�G�m����`�*��geI�jTO�a�0�:^���}h�/�u�9��aL�j۾7��|5)xw��:�< n���Xu�B3��e�b���GI6Tz=]��r���ğ�
�upvJ��1�� �*�tM�D���D-���ԡ���eb����t��������!8Om���H^���&7�薭1V3O?�	����XiJ���},N3B��Da��.n�m����Wn�,��u4���+ac-u|6��73�GQ�ʺ_K� Ϲ���J��R�)���<c�o��
=.��^Lj�"o'@�;���8��]�M;�E�78Al᲼�$�E�wA+� yټ�|j���qW�%d^���uS�m�^폝�q
�V	��]b��~K ;�j����%l�Ԙ+�t������J@��YD�:���V;��T"��a�~���m�)]�2}���@�{��`&�n�y����%д��뎶j�D)��,�0�c$�'��g|�m<�HM)�EaZ�Tv�8���,a�x�$���B�x�X���S�����>��� �##a@=A��͘��{�����6�ع:�a�PCKUY?l�E��%��׵1�c�XӇ]O�N�m����R�/m1�}:�������~�,?���,32M�l#褳A�]δ��ܩ��3���}ۇ���v�<�5�^ �����\c�dE���~�<��Q��K'�	��ޢ�����;j���t�!:�/u4���Ng�S�K�?�r�,R�5��c��(�p��+��[�c˛Z�ݵ�[9Ji��j$S^����P�HY��I�N.s;�2ٕA�X�E�$X���㸼��[Ψ6՚S�����+C���y�FG1E
,a��9:��h�����(
�/~
����fG��%�zY#S����a~�j8�8Z&��E�^0Yhe(�CƊ*;Uai�N��7x��|lzx�A�
`GԮ���%�E��X���H�S���S�|m�'�¶�`L�"�'�����!B� ���|�����LI��(�b�x���wtOwt�j��~�%�JY����r�՜��6�,�Й��T4�U�*-��{<-�˫sAC�t:�mX��Z��&Ɋ����5����=(� 7�U��8-�6/Wy3^4��wfM���yK��|�N|���g(��SJ
+}���f��0Mp?��TR�j�w�5\���r����C���ң���Z�?g�X��N�Բ�~��s�w<�g�)D�HXB?EL�.Ӄgn�E�����Y8�$vY>�ײRŐUU��~?�:UT�v2��珯�w}^�˹�\��H*�LͰ@�W@������� ��~�'�?.]�1D�\x(?�z��i�ŭ���0�G�]�.��i���"M~~�7i�S�s�#���w	������XY~k�k��t�����դ�*��D���/��9���i���GH�>�)�/|ό�p�g������	%0�I8��L�{%q����<x�`��:�E%��\�3���DӅ��)Y��a�%�t[:/]u+�� �z�H�5�n��=	��#xb�)�i��F�E�;qT�xE�����	b0m�5���9�F���,km�⣝j�Dv�u==�Y����b3�m�
є��:�ڿ����O�=���=�ߵ�I�[L#n���:�p��l��&(��f}�4Ϸt�#pj�;�I��*��L�R�m
Tᾊ\��qP=���̉��G�VXQ��E�M@l�$t�Q�\��M?+!N���Ԁ��9��;NA��JY��G�v���� i�U`��O$AԿ���C+���7w���XALo��	TݶY�h���R~���<���܉H'�.|���i�I�n���,>CL��c��AJ`NNj���Ʀ(�eƹi�D�d��֜&8x�U�ֳ�ekRC����n���{Q��˸�[�2�ѿI��.��2e�x�,�
$��Z�e���
�e��z�Gu��p�_�c4T;�����\J�0,ą���,���YU:�PfҾЙ9�V9qߜK!'���,��o�zN��B��DÒ��[��-�d����_��# i_��c]w�V�G^ �Q,�b(W��{�}fW�lC�L�p2[ιL%(�5q|0F����_���6 x���N�Z^�}�4gְ���q��UJ�I��4"zB���A���q�2��;�u���{�.����T��TQy�#�UL��/sc�y���t�l���@1~A�$��v�K���ܯt��;�8�oa�����|�s��Ǉ+n0�d���ykV~e�\�������NFk@�M���b��T��g����kk�2�q�&ʦ�'�u��Zc���?�-U��k�$H���ܬtX:�H���j���T˥�]�����2�I���o�ׯ�Gg |�z�������� )r��V�D��:I���ʆ':��(��Pwg���6
?8z!]�@'l�6�7��͜�a	�h�'&�s;��3K����Ba?�}�Dm�7�#aM�d{�!#��HC��@��JD������.�
��3QZ2���Eax8������䘖z�xy� ��
�~
��OH�)kv,��߻IR�7�T�����婖SY�m�^g�-݇󸣖�na	fͧ����R+��0
hI�̐ϩ���ǽC�]3�ʿ��/}�2��Cl�P�2�5:���e,J�@�]�b���B�o�a�n{���xT�)��c�6��v�2l4�A�
�
����H�}!`��� ���<B�U��̛΋*�mtBؐ�w�q	�%�o�-t:����_�ݾ���j#�VA�h�M���<�e��^� ��� ���	�Yp�E徱<��&�9���!}��1�]��}����Z2+��������?�c�oua���+U���[��y&}�ȶ�B�H���dϳ�=@u���fOE6��^\��h&��}�hp��W"��{��~�ЍE�W �K�
���o��K+��V�fwpx���*ry�(�+C�}�n����Ȝn���Ə0A-1�t���ϨF��lK�lR=9����S��hL�U%k�7�}�Rʼχ�nmvc�r����	⿸$e[����A�E3���lA�c���`����!�&T,{Z�,̔z���%�5�x��[�zw��T[^�C�p�޹L/��5��  ��<�瓉r'S��ң}&��ח4�Y�z�s-���4S��+�1c��l�Wǲ5F]���a�ǃz ]xd��ڴ���6M�_�bP� W�S��-:+�X�fu1��s�� jʻ?�L�k�����HrD�-{��<���A�4��� ���28�Uk,DPh�}�-����/�r��WCNؤ�ו��e����#8/��̇��),GR�E�4�*�x埾d�%'�~k�7����{w�gKl/�����kƋE�!p��H K��^���Ef�H W�3���i�B�&.ɭI�ܾG����yR'h�jc�����p la]Z:؟���җT��'��	6N="��}	�?������8R,��o�܌����k����&.�T�R��$��&]W�vQ�M��虫��,��خD�d�+�
�e�d���ߩA�V���z�
��F�*g� p��FU	���"L)p�0��Ji��Vg�[zz���'��4s����L<I�K ��>(v�p����MYŻ�[�u��S�8��A��D�-��b���C�,�q#k^K*�g�T� �=��cTeF� �랸Pdb�	��8>�^�
S@v��+u9��_�ӑ�/�q�F|�^�s���f����:~��B�;��lߛ��aѪ�J�V_7ʃfY_��5�8�S�V��5�E�e�zo�q�Ũ�Q��g�7I��� LW٥˙Lfc2��X�C�D�򉕰u�ʇ"��ح�I8�nka��R���3���M(��6���/�!Z7ٴ	���:�'�Z�N�8�)kjB�_-BAtN��(Og�k(1���uRa@��y����3����J���O��CJ�j�nD�"�!2��j�<<��lP�V2	��$��1C����6�|���:�$��R�L��PQϚcr�z��a�����M#�vGm�}�g����Yv��� ��w�%B��apg���Nz�����]��MW9d�o!�&ob���	� ���Z��T?R��HA�9OV\� oR�`�%��$����@��T��i�2�uMQcI`�h��_���E�WF��i}6?�q _Ym�S"��U�<G�2�KJ ��]�&���f(l�9 ҥ-�VO��d몂V�FB �,���?D���B��Ne��-�B\*i#�n�҃e%<ZH������[1�Cpߨ�H��neXf���,���a��0�y0J͹��*&-U�(��J@��{���Ӓ���=<`FQa�@"�r�f@��ґ��|j�r�d�p"�82rԬ�wޟ~���S�3n����p���OO���e��gݳP��~��nbŧ��k���#a� �5Hc{�ad��9����n��5N���TטsP�&�ﺄ�T�2'�`�k��x
h�tmeY�y�%�A=*Զ
{+T`"�K�D$�:�.�̂��Yߙ
����(P�މ�"~|U�_�E��ɺB��*��ӀH�`p9����g��^����{ް���F�/Ƃɡ�Vg�>����P��g.[�oޘ���Ͷ�
Ά��f]\;�α��)a�t�䩜��-%�=[�������ﲝbs�C3��f{&_��i�-����4O��ih�G��X7((�E�V#�>h����pP�%��X.�`W�B�@������2m�=@�rej]t�i����sI�7::V�N�8�VgL�������Gp]k��;��+K
X�p�ک ��0���t!��Ftӛ�^�5]�r";��Q�	
�<m���2�N WW9PM�Bw�Д
�����~8^���IY}�E)#k �j!7f�`�o�]���Mp�Wa�׶U1�Y>΢�lfuH�28��eܘ.}	����wb\"���ie�6������0���iQ��r��w4e����=G���Ц���pZ���"�8�Y�J�z����#�l�!�Q�*���گ��˴�����D���Z׎�2j�[`"+�?���I@�Zˮ���^��a8S�9�֡v]����		�x�z�!v$�'Zj�q
N����i�	�d����'������"�;�%IJ��5Wt�V0�+��$��-���ܨ{�_RXQ{�e��0�2=:��6qq;q�S�l�;_�D�i��e��(�1A�p&����_�4x�J83�$��vzv@�e��޺*i0����ƙ�bQk`o���Q�=#�lw����8qr����m���wr%���w�,s"�?�ƑZ�2v��a׿`�|d#���-G3�~��2�k�XZ�B{�r�"�!��CW��9-��x"y�,EI��i:��T��y�K�a@ڲ�5E�@O��e�v�3e�> sİ����.��e�V�㊥��O�#VݸĀW_�����p�n��j&r��O��"|�w0b��^�o�n�q�w��6�^�E&P���XB��ퟺ���NFe���#qe6׀��A����l��=�ڸ:�/@��d��L'�ͻ�4	�5���M��J���l^t�,ֺD9{+<���݌���k�r�G�Uv�d����S�6C��C!Q���l
��\�Ω�O6l@KFi��F����q[�kh���*��@�R�^��,	]W�	�޾qL���a����|�l��3�����~?(��
6��h!O׹JāzO�%se6ߪU�J�)�H��1�,�������T�#�N��2Uwf�Ȍ}��Ŗ��Nn�r��L��T�{	�P-v�D��'���{����}9��"+�un��Zl�p�o�J���|*�B���EƩ�Q�M��TTX��<��p$��0�۟��a(���+g"�����EU���2�]�u}�(B����!��B|����)<����m
?���t0vd"�/�}:JmV�����rA(����7`����9V!���X�?{���s�'��2u �.A�Dp�W�[q�7����]�8��(5�{u���H��ې!P��Κ'�׭O���3��Z�����_����J>GdFs�f�����ɮ]����Kzԩ�Lٛ]������G�z��{7�v�������*W�}F��/<����^������P#��XnO;���{(5�y],(��^0+��a��!��)���S���������ݢ: }4(=ن�;`�/�}	���p�)� Ȱ��s���F��ކ%<�9���m,�_��銦��'�]��ϸ�pkİP�|��!��"��/����0<p�����(tٯ1�7���� ��~*[�>�wR�p!^�$��v{�\�|�AM~EW,ȺPF���lמ���nj���J�~m4`E ��w�eI)�r|\��@�[��eh�W��?�8� `O˜��sH{��tA�I.�.2�������	&���k~��%�ə�{M�`�)
o_�i:�e~T�T���|\<�Ų�.G�(��~����-X�ò��� �P0�����U�P���1e@���W� �o�(�=�G�V ��������{wa_u�g!�7$�?��R#�m��$��n�W�p9�R઩i���݊�<[��cs�0N�MP�E���n�_d1�F�����ʄb���/����	?�s��6P�qٻ�9��u��.�J3@�����Z�~uܪ\�P�S��&Z�V%�^Չ]H�v1�E��WX#��_���7*�F,Rt�{S|Ec֮��^�w%?5��֯�»��[!�_�{<�Р#�l_���6R���!���з�P �֞q�fv�pf�C~,0kk<��Ѻ��
�
W������6j-�Aa3�ajmN;���z�nCGćj]�r�8�[�׍!G��&��kt�����RG��:z�?����W��W�UʃZ�) ��lpYp��~J��gbk�!&w�x�-~g���@�L�GB*�ҝwli��V�y2,��p���V����/��������\5�~�9 �ÆD�>CşX���k①_aO�T��݋xA��D(h�3�Cw�%�q�_��>�W�0�DP�S���4�K|̸hc>9Ik?�Ŏ�J���_��`�NT�K�`����G�I������2(7G�J��ЇD���+c��_dN�Fގ#��߸-�w���.l$�(X!4��q��-1�'��9�h��ֽ��u_�~��f�?W��@��t�c�t������I9��)P4������C�^v��dn0��q���&{aАY�`!Jc�)��ھ�K�ۖ�y~�w�����*Zǀ��G,���T֞�����s�6�����E�T���#�η�����;pA�b=.���ʋ�#���X,�*O�����0;��}`*�dN��V9�����
N>��+��JQ�7 z�kS���*�c姼�g2b IxC5�S�;1��S
��Kт.��\y�1�ҩ�g���:Tf ��JI��ke.�T<<m�Ɋ�c���֕<&���PT���[�n�\�촇�������v����(��+=�#�<}D��^BT�R�5R�0o$��->u(�"�I�C�F��]����{��D�?�=z�~h��H1���8(u.���Y�7��� e�V�L\*�RH�D��0�~��8%Cg�F��,��Y=���!Rk�� >I]�*- L}��J�W`��פ�)pN[pl5���Ɍ�@c�a47�����ƱG�.��!*�A�d�g����
�0��F��27SGoO-��PH�$]���pe5]\@1^����JF��j8���>�	��*TS�1�
V�"4|�F5(��r�`���zO�r�я�ʧ鉑d����Bsc_�sl^��	�D;�cK�`N�fp�\�w���k��qE_&';T6��><�k�&���Bړ(˖rxgF���J����dZ�$Եo�/�QMx�0C���Q��T3(0Ud���wt��۶��ei�z�-������R,�i�Y�_^�f�jr��W{ۯ��5~/�#�\|И���+BJ�k����w��H[�J�-�FV�����,5!f��O�J����� �D�����k�q�9�5�;$�iY�Y*��dj��w�;njÞK�	���c3�^�J9��Mz�H�1�����d���02��٘��6YR+�}���^9���< �rv&Prf:�}��=HI:���@�K�dI^A=�	���?��/�s&��w'@�Rԏo2����a���.`\汯�>��=��S��`�Y� ���(�Ѳ��uT�4&�6�a���Ҹ�9�O��enN����b�'�+L�ڏމ�]��/	�$�3�]C���~��������G�HF�l�A���2[�5��L���_<)#k� 
��2T7^7�:A�8�O���VN�	-hbW�n� (��R��-`/ɇY�4��]?��d�ڥ�f�p�=�s�N �����5��CC��v��Y�w���?s���N��"g3�6 \@I!�ݢ�a�̃3����
WJ�h��FD*�Z9_�Jv�#�](�@y4e>�s(qa�4��o+��
|�p,a���!=��+�-
ĉ:z^�ĕ4����mHkRlh��'e7���TT�.�0����g|k����{@�����x.�$����X�a2#�dD��CK\r/2����;QM�+v��b���<����6�Ih�U[R�]�y&;*"�S�q�4�G lh�uZN�� ���]D�2|n3j$	W�`(3��W�M�l�m�=��w��/0n���9�����;� �)r-U:�5d���9�#Ɵ���ԷR���Q���&�������t(y	X
����֪�D��v���9����۸1,�q=�0G������Y{����_ib�9�C�\'�r�=�Y�X�=c�5C����K�6H~���'�٥KJo�݀V�^`+�
�ͽ�M]t��W�$����TF�[~CM�G3�,���a��9���'���6�BY�x4��!-���%��zo6"������"XӜ��m#uGJ];*Ŧ?��3��� !�-��ܞV˫����#�Cq��T����4W Q�,`�3���4��t��7v����TDQ]A0a���ysݣA��C�e�j�l)8�I���^���J}*��^՟���mNqn���}�Y򧉦k܂u����["[�4�>ޖW+Ӱj-/��16Y���Y.z$��[�� ����s����F;2��V=�6�K��v<^�5D%�`��S���8�nY3Ƞ���
96��v���/��R��}��Пe����D\֥�m��-1�4�5j[@�&s\h�y�M(e�
s�t��>Y�����MF��pV�v��y�G��gs�v0b!ٜH ����|���B��U�*IQ�鷽N��6��]V_�j�Ty}l�9�P?D0u��02���D|����!�Ӏ�ɇ�f������� L��!��}S0e�-������