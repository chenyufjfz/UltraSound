��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>Q�y�`�}н龓I�����>g������w�O�������x�d,p�ܞVt�}�񺮻�G���-)?������"�c���x��B���_"2$[��m�8��H���`�/&���
{�90n��2@����4���������#�aOQ%�q�t��6�����=���R�j�7���fqCc𞴧���c̿����#4^d�X�*�%7�2�P4G�(��uI$����(�=�r�©P���	�/��-(_�65~i�ԼA"'�(S���-�]`�~�/�|ea����TP�h�㏂\&p�y��V��A���jpDe΄����c&(_Q�8�z��t�`K��N���%�zC�z�$E&gJ�y�?Ҋ-�b��JH����t*ry'��0�H,����'+g9T��{{�S�+ ��� ���3�����p���e��P��P�I�{|Ҽ����Z:4�e�@\ ;04�j.s�N
�,u�ƌk̟���/
���������Uћ�[�K=���HC d��j�[KW��m7��&�*cI?�����:[����ޯ��KL+��qV�4� doXC�8'�9�TXs�!�4-b;��?�g�5��>�s~   (*�\r ��6�����~`.�X>>{�Uz�1��"���<�7��qU)\y�J���J�K���B��?I��j���LZ��)��3m�țB��.�s)����/˟g���wd.��0L�VV��<L��vԑ1GC�L�������3�?�	�4��<k;A�:ѤT��L�
ܠ-���[�f���d��-?�kj<@[��ܧ2����J�"��!������?b��o�أNv��-�xŏ�␢,�t�D�T���vw��9�<�="9�Эީw���f5���Na����%DXL,:����MN�ȧנ���z�·`�:�`�A�+y�:]���;#�p���Z��B��W�Z�eiy�[��w�������[E�)'i]l{�='␈��|&�K��oJ>?�/�>�f���U�N���S'ܭ����Z���s�w���	��v�qn",Z�5�y�hi�!���IjQ�7e���+n�u�4�D�`�$3�!�J+YM�]tΤAT�qS'*�+��� �k\4I�hP��x��!)��=x��M��,Zk������)U�hy�-��e����@+|�Y��Lr�|���Y7۽Pޥ��R��ZS�}�W�^�a�����Yz�ڡm���_9��<�p��A��,b��F$��w�:��E��j�&�a)��m(U�kFD��)8�^u6E�^pI�&�>�Ĝ�[�*��%k^�A~`���Y�p��.�k�����`�]I7ð)<Gyl3ZN�)W{!�� � ����.�Y5�ʅ�KxIJCJ䂨�kQ?��X/{He=^5�u�bn��D�dV�p���S�QX���:��;�=��ft���z=hd:����{p�x�ͨ_�()R�.Qc����/��4�9���N���*�$��}V:g�wx�M�c�/RhZ~��~�6[��ـC�v3+ɴ�4�.$I�4ϒE��,nX!�TS�?��`��[N�WZ�8��!��x��T�14�:Hk?�P^�_��tJ���ݓ1��4װ��/v�q�ȁt����;�#n/�<Jʄ��_��#��ᕲ�U<rv@�|#��buы�+���NVe�������P��3�^RS�z�irTN�4��Sq	������k#)������L[�4g���S܀;b��#Ac�?�V��b��L�����x�NԞ�g;��F����l�7���#x���>�_k[����J\ѐ��G�`϶�ɝi���!r%_����,fX$��sȴ1��b�����Ug��p�3�g��I�z7_m"k�PL�����h������&�$�d���g�B~@��MF����h|�����9JR �ֳ�S�uq-�-jO�CA�� 2�9�E�"��@%ޘ�cCkdI�"lA3���eJ��h ��T�A��0���3+���"�x�	�?
��U���9�ٮ���p�:��|ndQ�G7w!��+���JQ�M��S��{j�1��q9c	��IړxyGE�f@)��W@1w�V�`+d3b��-"~G̓�L���g0w���Q�q�촧IPF�_�φ�N�i=rb��g�/�6�c�?֞��Z�bS���_����� ��07�N�#���V�Q�H�s���}K�M�(�TY�ذ
l�tdʢ�~����Ke?�q��U6o~^�94�ti�l�R�~��=��~w�
�+-�H	=�	��Kj7���-��P%;�F�DArT��
�#SM��P��Ev5+�w�g�횬q��R��rb0�g��D8��6����O$\~�����+T}l�4$Q��0ʅ=!��x��:��]�F/a�M������y��kX82����.�?LgԖ�'�>ی-�"h���3Լ:�)�˥�As��8��+r.��Q &��K+'��P��p�pO?8Z��Ǉ�i�"E��L�XxX<U�I�k�p�2ᓬI�uBߵ�u�K8 G%O2fE-0y+�E��n��Y���늶�~=k@Xeˡ�{�S� �J�yV�%���xL�̶^%wx��U������t�N��	�����z���/��?l���-��;�>���z�P�>���0�D���tW�\�����Q���a�X̃�l��?��+Vng,xI)�6-�ֻk�=�s_Ix|3V	�5Fm�8`���\��]'c����8��O�\'-6m�E�pO��8-��B5;�rʼ���ϭ���T��hx'��<-ta�0ŀ��M�(UHe?� g��R;��(}ZIϏ�^
�2�.:�jG�y7\������ɐ�ȱ�z7
��%��ύù�H,u@XmJ`�f���bZ3����E�?\�E�4���0�-���#f�:v�� Q\�˘d�h����S�0ę���9� ��*b4��v�3?��jp����]1�;����>�Sb:�;i��-��O��x�Y�ZF�k'�:!�m��8�?�k�/ h�����(��!/6k��K+^�����ڠ5�#dą��v)���^Չj��|e��H}��>��c���Q�8`v$7cwg��W_�	��?�������T�����a�J�F�5xe6�%HX4^
2�ါ��?n��o��K�K��C��2�d[6@�Ұ�(n�-@���)3ѝ�v�[�tɏ}o/���<ak��'�%G��ǒy���^`�"�脘��U���}'&J�qq_=��'�t*;��|q
&�E�'"�Jb�υ��΂�!�(�pK	�tҹ��ȣ	dk�-�sڣ�)Yn���u�1�@��[��i �J�-Z�ӧ��Q%=<��8?IZD.��c ���O��+�Ӣ���l�=�$���.�n^�-Y�?�
�ͩ��Du�`Z!3���MU�7��W����?��k���'�D犯wjR��lCBȿ,��N-���V��l{���lW|��5���0<��lx��zB�<����\1�
��$�#M�jw���VR�4�2���_����3A��M����ڿ�"�|%�*��z�c�)����ݵt)�v��Q��x�$��O�s/����H���r%�#�����X�D^�n�>\̲ mx� �q�"ME�!S�H��.�`��*�	gw��+���H৬���Οv��X�~\�<��?�
Qi#��V\c�ˉ�����ݑ�O�H�q��Xﰤ&7���]V~�ʲ��qU$Ѿ@��F����7*U�%�?�"�l��o�h�2�K����HW5�/pt��ϼnD1�hK7�V/g=k�]��	��$��
�l)�p�猎x�^��a<=����D�+��9l���1c����2p�K4Ŏ�ؖ��[qF�������}�?ݡ𹶗 Z'k���A�EY�R����q�Y��!�-�3q �Z�]�0���n~��Q��'�0V0؄��JcfJ� ��݄K�����{5���+���BR���i-��x�lM��0���:l���5� �c��̚������������i�QU2�.o�_�;7��ʀN��_��D/�/~�ׅ�RM���g���[d&��+Vk��"��G�cB�`�����m ��`驮&ԞIgAǤ�
.\sN*�i���3
0�ޔ�������K8�R��@�� ���~��e���23���8�,ǡ�x�@��:���5Q��h�ɣP0�K'E�υl��,�s��G.~����87�?~�Pgx��q��"g���1G
���y!yi��넺�mjڜF��d�m�F�b\�m̧|N�*��������]>0Δ�ӤY�2&�����9�n���(,��}$��jBl��΀Y�($1e���b@��!%�Ϡ5�b�BI�gM�� S�˱�g�n H��A��SE�{k�z�1*�V�����b�C���"��RK�P�ޡ��{����n�ME���rC�I&?�A^(�X���Z.m�!��:��[��h5�_u�)�/,җ#���U�J��:��(��&�dͅ�m>���6���65;����CW�-�q�l�3�y�YV�%d�_�4�kH��6�ٍ�g��k֏�r硅Wi�	q3"z�_F�D���8�L�����Յ���0�mT�D%xgI�7�p�,�ru�����r� v��V?�R,�Y���a!-N@G,��f��9�s������_��
�0KZ�����Dx���[f��� 
��WZ2�l�&8~�O٘)ԪI�*�A"�c)��d����� ����XC�� 7,zX���;�T�!'�R�%�6|Y���YJ� k���W�����@5<��RE ��	�Ȑ28(=���^s�P� �I��˨d^:���[�_�La��p�����Uqp7��[���pA� �sI�yh��?�c`�Y�=Q�F��n�/^w�EFn��R��{L%j�k(ّZ�?�:���nG�1�r&�dL�ig�zR��`m�,UeR�ٜ�0��"h�V�RS�u]�[i�dq:������iPs{F ��Sc<P-�����&܃��[Pc|�B� 7�:���;v�:L	���xdΒ�
B�����_�YH"�{bV�4��9�M6Ks��������^3r�E�}��}�t=��r�Ł#xvɭ�a��3�����3�=L�쬕��q�F9KDx�&z}�@�ie��|
��z�D`j��]9cd0Ckd�@ �b�ٷ�2)�8�	�dU������f�b\ǵ�jF��v�_��� �p�+��A�TS�ϼ�(�K���J漋��*�.�R�|�HJ{��<����эx~k0��J�e��3�8����6�J�M�v+���2�W����8�Q�I�d���?�OP��Hk��}(wY��O2jK�;�u\�w�H�>�:o)�z�j��kP��q�*�+��SI�l��\�;�� ��$/�. 8f/k!�[)#q��x���	��:
�r>L`� �E�\�,���x��n�7*�F��wv�L��*1����0��{�t��=^�$�k�0�r!���'�g%��\f���}߇\����_�"�#���q�%�
��"!b�e<�2���
H-H�'s��9�z�؆����I�+�wK��jڗBz���L�]��<|���Yߍ:&��DD� ����_Ѹ�����o���dhk�|^�Vޣ�ш�HW@�"NU��H""�L���p���[X^֛��'�rY�\M����!�3�l���Y�N��]	f2���!��+��5���T�D�?�Ͼ4E=�3����^��-e��8[j�GuDj�1$&�Aq'e�=��!tW��Im�J�k�{,)����%����q���ch\r�F܊�ᠣ7����͑FL>^��_�P;��t�@2�a�1��T=�hT�e�'1�$5��;%w0����`5��{��H��<-f� 	�\w�n}+��Y���d �^�cši�;����j�YU��/`�9G�}u� ��@��n��������ǩc�zG��m���JN�/C������cF�T����T��u�
;�s�Lԕf1�%�r� T�w��%k��P63}��Rzt�.�<�I~� ��٥��z.%gc����>v�S07x�MEl�^�;��E�ԟ����{cU�4ZB4�D%�n�Eɯ3�g	Np�Ţk3]ߦ$���=��I������tM��*e��^�m4�+���{�aX\����+PVAu��"f��昪7qP�V9Z�*]��m��.++��"�y��$����jK�J�D�W�^��`$�vd�n.���G�#��m�Q���
�#ye�w�%���-�&���M{i����;����2/f�@KtG��	���!m,�}R����E�,��0���i��A���i,�Q@Nec�^�}��4[��Ay�KuZ��H�#U+a�nB�7�.�Yx���t8���9�H�J��2ϾF&��Kl���`L�Y� ܊dHe�/�kR�T�Bz؆%p���v$�j�'��Y�?)^N~)~���$[,"�C�V�v�c��*��W��tQ�s��]�ǖ(ѝ�)�:�nY�g�S�p#M��_��|�/?>��ŽV�v��Bgp�H/��g"��Ԓ��7[����9�rݓ��U���S�tѕ~ǳ/!������k�����Ek�ii���~;q��B��5oDS3�Rp���y�3�3�PL밶�g]8&Cԑ�#��}:H0��[IVic�T"�|$��&<˗���8z��E���8�Ҭ!NlĎԩ_���et��ү��F#z��+�@&e��9��tjP2���P2�� 7�z�Te5��Џ6����*���s�Z|ɀRVdl�̨^�Я}S,�Rj��n�2�����9�?O���,T���?_� pͥd��8A���n�ƕ�bXAG��m�+��g��;��̎���:�T�k����R)zXGN���@$�Oحcz��������Fn����K���L=I����|�x�\Bi�3~��ԡ�]��T@� jƚ�r�N65���o���b�KMe@l���6�&�Ј�p������KY5�Kp���?��y�ZT��¨�c͵Ė����F$�KLF�a�fVǤ�zD:<}{em������Wn[O�c��+�@�[���,��� ��F�˳ozeD�9�r� /!Ϥ���Z�YP�xܸ5�.�.Ę�U,ߛ)'ˏ��W�u��J���ޏ,���Z-V����HC"z�gf$��qOL6m�[B�X�J֙#���bF���7�������E �p��3� }��U�qz-�����/���[����'�k��l($'���vպ/��1����-.�l@r��w��1�߃+D~���u����]����u�[��W�FL�c�:���OB��{�S�f�|,���v�#ł.k� 7
�a�,2�KX$�K��XP\�H���AC�҆�3M�2BkQ҃�:+q2F�r���m�B9+����
��p��m�ة�[1P��ۢ�hp�>};V4ءX� h����%{N�GFF_���f��������v�"��:��좖%,>�A�>��E���6��f���������H���f�c��t,���O���E6�ڝDԺo��T1w�O}6���T�7*��cQz�Z��N�;�Wu%�JI��^�{�ir��(���ߝ���y-D{�${��q�om����E���Ĕ�r��s1򖤫�'�{��n�L]��:��
��<�ڽ�|��d�`�%�R������W+���k��{�M���W~�0�W_��D^��&���8<�8��S��@ȦU'4+e���� �8>�`R����(��G�.:�fE�RUC{�{G��6�'��]�%d����qzHG�H��{8O��i��B�B��������9q�~m��X����8�3Aah�����4��%X�2�rs��"Cm�>�,~��,�|a����]�<]�[�٭�L�x�7oϬ�v���睠�r�6Nu pSv��U�7�}��� ?��)��#��Qb��ŷ��+��� ��H-�HF��l�F3�������$^�_9��~'ƶ��K�R�5�B�e�V��k�����t~mo�|�v�X�~���M�=�w��=��!��csvDsH����e����ׂ$����"�$/�I�a�ZT��	l��� �_�+ j0�^o"�`����\g�w�)0�n�*ɪ	a���5��Nu�a���T����v����_�о�Z�7�1]��N����Ə~�uӼӳ��̮��� ;�]w+��_��R[&ǈ����� �ru��-le�5�����3D�L'�/�+u���i)��H�`�����YIp	��_uF�A��9z���H�5�O������d�6��u3ݛ�jC�De�����\�;w��L��X��8�4��/YD��J�
xK���S�@^V6n	��7�z���d�U$RC�_��G�ko ��O�� X�������d�_�	�)L]D�h�K0�̛ܤ�WI�^���E��n��OE[[�W>���	 *I:�|y����1PE���R�V�[`7�P���$�]�Kn��P@��Y�\���#��^�"_����rr�鏱P~d�p�1�^t�X�s���A�cT�.���N`(�>C�<!`nYs���a��b�����*W/C�}���Y�{'X���#\�z��;�����ٖ�= 9��R��I��n�����e�sL,��N-���a��,��������M}�2��;�ßm�������gHq>��!��c�~I���yAExG��2O��3���E�C��V�^8��
O�a$W�n���n�f,�ZO�)�0�3��(�q<Nx@E�A��d�P�볶P��ݶ�:n���Q)�-��/[I�i��.�?���E�T�l����Y}�`�)�3m�uZ]�Qp~Mv��Ͳ�ż��܊����{�k�YK�刜$�_�)�Xq��6^�٢��A`n`��P�*�j����+,�"L������fKDP�� ���%����Ek;Spt�K�C�uR"	=�kͶɌq3K�p�*�����& �'��;j,���$^�0>�Nz��^��R�S��ƈk��MAI���覺�_��R�/��*L�nd����t���j]�7}����������&S/�XUNr+e��1���GŦN�q�R�f��i�xN���o�Ft�=�IЀs��߶���z���~�[Y7��Vv&�jHt͙KV�y�6��@��CE=5�(�U Ǳ_R�\�d�6�����!gك|c��%�O�hz�E��2�ud�Cm8�/����~d���U��?9/ʍ5��̈t��O��[�X/�d�ܬ��zMd)8��{�V���!�[�l������O��¶��v��Y;M�tQ�A�G���󁺾�lsЯ��"�}n؊y�]�$����>BsRye��8�Q-&2p�.����2���Ѳ��oc���:w�>��i �,,���"�zOe4�tgK�0wj�mA,���.������ƥ���Qvd���4�_x�Ω8*��\�$����2� ^{�P[�nnˎ%�N�E�$�f?Y�KC�5#�V�g;�ns�/��R��9+�NRM]tkU�K�e)=�[fWU6�؂f ��������U�'�s��%����yoK�8!M@���+�q�J��rΤ�y�h�:�/%tj؜���g��XZ�+�Dd_܄����H��5F��!TwJl,�j���e�=�R��1�c,;��T+e���"-c=�^�w�������ճ��cʇ�7�&�T�&�a��=Sa�C�w!�ʺ�q�[��J�x�--�Ú�p͌mٲ��}���K��6�n+JQY�j򥏁�P_�M����X��ŏ�7�%��7�>}��%��K��&���o�v�@l"o���*��g��pq"���n�0Ojҁ.��Z�mtYm�6��o"�^+U�ׅ�Zl�HI�"�w�\���U)L"�5�����Ak����(V�����.�SI!]фHex*2x�b�Jx���s�wD��հ�E}�����X�+{��׭[������^�/�s����P3G,�x^>����O�Dc����c��\Π�����Dq�Q���KQ�� ��	DѯJ#�ʯ��Ht���KF��)�2U9���"l��]aR�a�P�d�$��G߂��˩A� ��E��!�������PG~p;��u]F[`&b>�J�I���X�Ӣ�m����H�+��ˋ���8�`�?,��4׌S{Xi6Q�+w*�YK��؉I�AS�xhC4Ԃ��J�&��g}B����wfѫQCyL��d���sOŻa�A0��n�'�����L��i֜���4\��Z\X��q�Ĳ5��?tRAͦ�4-˓9�vј�ee�{�1�P��r�%�~�n��ģ
+,uH�_��������u9�3�
N��Br�Gި:�D���@WN%COR���,�#�i�&�V���y��#ξpM�r�Z��~�J|��6�������,Nղ��ŉ>��x�YF�C��x'�
���)�x��`]�˟[}h�_F0��ucw�1�]<�zI����p�r�n���T���B;��!+ui/c4�����/%�	M�D�K���ޡۤ��[ߕ}Ĥ�е(�9S���+�%�Ws<�C�/�?F�K�����ӭo������n9��vA��q�c*���3��
���>IP�e4"����j�� 6�l�id��B]ֱ�-,=Y�UcJ�.9��60��gc��YX� 3�s����4B�8�l#�Y�
�g���2�X��C��Al�'/�uM\���1��΁]G�ꓵ'�ۦ�#K����0�Ш��V��/y�}���<@����&��+���:+��u�� ~��`�(�-�0�b�\+ղv��N���Ǟ�&�w �O�g��D��|�-�K�$<3a^��c?ie�D�q