library verilog;
use verilog.vl_types.all;
entity udp_complete is
    generic(
        ARP_CACHE_ADDR_WIDTH: integer := 9;
        ARP_REQUEST_RETRY_COUNT: integer := 4;
        ARP_REQUEST_RETRY_INTERVAL: integer := 250000000;
        ARP_REQUEST_TIMEOUT: integer := 1000000000;
        UDP_CHECKSUM_GEN_ENABLE: integer := 1;
        UDP_CHECKSUM_PAYLOAD_FIFO_ADDR_WIDTH: integer := 11;
        UDP_CHECKSUM_HEADER_FIFO_ADDR_WIDTH: integer := 3
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        s_eth_hdr_valid : in     vl_logic;
        s_eth_hdr_ready : out    vl_logic;
        s_eth_dest_mac  : in     vl_logic_vector(47 downto 0);
        s_eth_src_mac   : in     vl_logic_vector(47 downto 0);
        s_eth_type      : in     vl_logic_vector(15 downto 0);
        s_eth_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        s_eth_payload_axis_tvalid: in     vl_logic;
        s_eth_payload_axis_tready: out    vl_logic;
        s_eth_payload_axis_tlast: in     vl_logic;
        s_eth_payload_axis_tuser: in     vl_logic;
        m_eth_hdr_valid : out    vl_logic;
        m_eth_hdr_ready : in     vl_logic;
        m_eth_dest_mac  : out    vl_logic_vector(47 downto 0);
        m_eth_src_mac   : out    vl_logic_vector(47 downto 0);
        m_eth_type      : out    vl_logic_vector(15 downto 0);
        m_eth_payload_axis_tdata: out    vl_logic_vector(7 downto 0);
        m_eth_payload_axis_tvalid: out    vl_logic;
        m_eth_payload_axis_tready: in     vl_logic;
        m_eth_payload_axis_tlast: out    vl_logic;
        m_eth_payload_axis_tuser: out    vl_logic;
        s_ip_hdr_valid  : in     vl_logic;
        s_ip_hdr_ready  : out    vl_logic;
        s_ip_dscp       : in     vl_logic_vector(5 downto 0);
        s_ip_ecn        : in     vl_logic_vector(1 downto 0);
        s_ip_length     : in     vl_logic_vector(15 downto 0);
        s_ip_ttl        : in     vl_logic_vector(7 downto 0);
        s_ip_protocol   : in     vl_logic_vector(7 downto 0);
        s_ip_source_ip  : in     vl_logic_vector(31 downto 0);
        s_ip_dest_ip    : in     vl_logic_vector(31 downto 0);
        s_ip_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        s_ip_payload_axis_tvalid: in     vl_logic;
        s_ip_payload_axis_tready: out    vl_logic;
        s_ip_payload_axis_tlast: in     vl_logic;
        s_ip_payload_axis_tuser: in     vl_logic;
        m_ip_hdr_valid  : out    vl_logic;
        m_ip_hdr_ready  : in     vl_logic;
        m_ip_eth_dest_mac: out    vl_logic_vector(47 downto 0);
        m_ip_eth_src_mac: out    vl_logic_vector(47 downto 0);
        m_ip_eth_type   : out    vl_logic_vector(15 downto 0);
        m_ip_version    : out    vl_logic_vector(3 downto 0);
        m_ip_ihl        : out    vl_logic_vector(3 downto 0);
        m_ip_dscp       : out    vl_logic_vector(5 downto 0);
        m_ip_ecn        : out    vl_logic_vector(1 downto 0);
        m_ip_length     : out    vl_logic_vector(15 downto 0);
        m_ip_identification: out    vl_logic_vector(15 downto 0);
        m_ip_flags      : out    vl_logic_vector(2 downto 0);
        m_ip_fragment_offset: out    vl_logic_vector(12 downto 0);
        m_ip_ttl        : out    vl_logic_vector(7 downto 0);
        m_ip_protocol   : out    vl_logic_vector(7 downto 0);
        m_ip_header_checksum: out    vl_logic_vector(15 downto 0);
        m_ip_source_ip  : out    vl_logic_vector(31 downto 0);
        m_ip_dest_ip    : out    vl_logic_vector(31 downto 0);
        m_ip_payload_axis_tdata: out    vl_logic_vector(7 downto 0);
        m_ip_payload_axis_tvalid: out    vl_logic;
        m_ip_payload_axis_tready: in     vl_logic;
        m_ip_payload_axis_tlast: out    vl_logic;
        m_ip_payload_axis_tuser: out    vl_logic;
        s_udp_hdr_valid : in     vl_logic;
        s_udp_hdr_ready : out    vl_logic;
        s_udp_ip_dscp   : in     vl_logic_vector(5 downto 0);
        s_udp_ip_ecn    : in     vl_logic_vector(1 downto 0);
        s_udp_ip_ttl    : in     vl_logic_vector(7 downto 0);
        s_udp_ip_source_ip: in     vl_logic_vector(31 downto 0);
        s_udp_ip_dest_ip: in     vl_logic_vector(31 downto 0);
        s_udp_source_port: in     vl_logic_vector(15 downto 0);
        s_udp_dest_port : in     vl_logic_vector(15 downto 0);
        s_udp_length    : in     vl_logic_vector(15 downto 0);
        s_udp_checksum  : in     vl_logic_vector(15 downto 0);
        s_udp_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        s_udp_payload_axis_tvalid: in     vl_logic;
        s_udp_payload_axis_tready: out    vl_logic;
        s_udp_payload_axis_tlast: in     vl_logic;
        s_udp_payload_axis_tuser: in     vl_logic;
        m_udp_hdr_valid : out    vl_logic;
        m_udp_hdr_ready : in     vl_logic;
        m_udp_eth_dest_mac: out    vl_logic_vector(47 downto 0);
        m_udp_eth_src_mac: out    vl_logic_vector(47 downto 0);
        m_udp_eth_type  : out    vl_logic_vector(15 downto 0);
        m_udp_ip_version: out    vl_logic_vector(3 downto 0);
        m_udp_ip_ihl    : out    vl_logic_vector(3 downto 0);
        m_udp_ip_dscp   : out    vl_logic_vector(5 downto 0);
        m_udp_ip_ecn    : out    vl_logic_vector(1 downto 0);
        m_udp_ip_length : out    vl_logic_vector(15 downto 0);
        m_udp_ip_identification: out    vl_logic_vector(15 downto 0);
        m_udp_ip_flags  : out    vl_logic_vector(2 downto 0);
        m_udp_ip_fragment_offset: out    vl_logic_vector(12 downto 0);
        m_udp_ip_ttl    : out    vl_logic_vector(7 downto 0);
        m_udp_ip_protocol: out    vl_logic_vector(7 downto 0);
        m_udp_ip_header_checksum: out    vl_logic_vector(15 downto 0);
        m_udp_ip_source_ip: out    vl_logic_vector(31 downto 0);
        m_udp_ip_dest_ip: out    vl_logic_vector(31 downto 0);
        m_udp_source_port: out    vl_logic_vector(15 downto 0);
        m_udp_dest_port : out    vl_logic_vector(15 downto 0);
        m_udp_length    : out    vl_logic_vector(15 downto 0);
        m_udp_checksum  : out    vl_logic_vector(15 downto 0);
        m_udp_payload_axis_tdata: out    vl_logic_vector(7 downto 0);
        m_udp_payload_axis_tvalid: out    vl_logic;
        m_udp_payload_axis_tready: in     vl_logic;
        m_udp_payload_axis_tlast: out    vl_logic;
        m_udp_payload_axis_tuser: out    vl_logic;
        ip_rx_busy      : out    vl_logic;
        ip_tx_busy      : out    vl_logic;
        udp_rx_busy     : out    vl_logic;
        udp_tx_busy     : out    vl_logic;
        ip_rx_error_header_early_termination: out    vl_logic;
        ip_rx_error_payload_early_termination: out    vl_logic;
        ip_rx_error_invalid_header: out    vl_logic;
        ip_rx_error_invalid_checksum: out    vl_logic;
        ip_tx_error_payload_early_termination: out    vl_logic;
        ip_tx_error_arp_failed: out    vl_logic;
        udp_rx_error_header_early_termination: out    vl_logic;
        udp_rx_error_payload_early_termination: out    vl_logic;
        udp_tx_error_payload_early_termination: out    vl_logic;
        local_mac       : in     vl_logic_vector(47 downto 0);
        local_ip        : in     vl_logic_vector(31 downto 0);
        gateway_ip      : in     vl_logic_vector(31 downto 0);
        subnet_mask     : in     vl_logic_vector(31 downto 0);
        clear_arp_cache : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ARP_CACHE_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ARP_REQUEST_RETRY_COUNT : constant is 1;
    attribute mti_svvh_generic_type of ARP_REQUEST_RETRY_INTERVAL : constant is 1;
    attribute mti_svvh_generic_type of ARP_REQUEST_TIMEOUT : constant is 1;
    attribute mti_svvh_generic_type of UDP_CHECKSUM_GEN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of UDP_CHECKSUM_PAYLOAD_FIFO_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of UDP_CHECKSUM_HEADER_FIFO_ADDR_WIDTH : constant is 1;
end udp_complete;
