library verilog;
use verilog.vl_types.all;
entity controller is
    generic(
        SIMULATION      : integer := 0;
        AW              : integer := 10;
        DAC_CHANNEL     : integer := 3;
        ADC_CHANNEL     : integer := 3;
        MIX_NUM         : integer := 3;
        FREQ_NUM        : integer := 2;
        COMMAND_PACKET_TYPE: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        sita_w          : integer := 16
    );
    port(
        clk             : in     vl_logic;
        clk_2           : in     vl_logic;
        rst             : in     vl_logic;
        trigger_exec    : in     vl_logic;
        ctrl_in_udp_hdr_valid: in     vl_logic;
        ctrl_in_udp_hdr_ready: out    vl_logic;
        ctrl_in_ip_fragment_offset: in     vl_logic_vector(12 downto 0);
        ctrl_in_ip_source_ip: in     vl_logic_vector(31 downto 0);
        ctrl_in_ip_dest_ip: in     vl_logic_vector(31 downto 0);
        ctrl_in_udp_source_port: in     vl_logic_vector(15 downto 0);
        ctrl_in_udp_dest_port: in     vl_logic_vector(15 downto 0);
        ctrl_in_udp_length: in     vl_logic_vector(15 downto 0);
        ctrl_in_udp_payload_axis_tdata: in     vl_logic_vector(7 downto 0);
        ctrl_in_udp_payload_axis_tvalid: in     vl_logic;
        ctrl_in_udp_payload_axis_tready: out    vl_logic;
        ctrl_in_udp_payload_axis_tlast: in     vl_logic;
        ctrl_in_udp_err : in     vl_logic;
        ctrl_out_udp_hdr_valid: out    vl_logic;
        ctrl_out_udp_hdr_ready: in     vl_logic;
        ctrl_out_ip_dest_ip: out    vl_logic_vector(31 downto 0);
        ctrl_out_udp_source_port: out    vl_logic_vector(15 downto 0);
        ctrl_out_udp_dest_port: out    vl_logic_vector(15 downto 0);
        ctrl_out_udp_length: out    vl_logic_vector(15 downto 0);
        ctrl_out_udp_payload_axis_tdata: out    vl_logic_vector(7 downto 0);
        ctrl_out_udp_payload_axis_tvalid: out    vl_logic;
        ctrl_out_udp_payload_axis_tready: in     vl_logic;
        ctrl_out_udp_payload_axis_tlast: out    vl_logic;
        local_ip        : in     vl_logic_vector(31 downto 0);
        pcm_udp_tx_left : in     vl_logic_vector(23 downto 0);
        pcm_udp_tx_start: out    vl_logic;
        pcm_udp_tx_total: out    vl_logic_vector(23 downto 0);
        pcm_udp_tx_th   : out    vl_logic_vector(9 downto 0);
        pcm_udp_channel_choose: out    vl_logic_vector(7 downto 0);
        pcm_udp_capture_sep: out    vl_logic_vector(7 downto 0);
        pcm_udp_remote_ip: out    vl_logic_vector(31 downto 0);
        pcm_udp_remote_port: out    vl_logic_vector(15 downto 0);
        pcm_udp_source_port: out    vl_logic_vector(15 downto 0);
        dac_cos_sita    : out    vl_logic_vector;
        dac_sin_sita    : out    vl_logic_vector;
        dac_choose      : out    vl_logic_vector;
        dac_err_clr     : out    vl_logic_vector;
        dac_err         : in     vl_logic_vector;
        ch_gain_sel     : out    vl_logic_vector(2 downto 0);
        ch_gain_da      : out    vl_logic_vector(11 downto 0);
        ch_gain_wr      : out    vl_logic;
        ch_gain_clr     : out    vl_logic;
        ch_gain_gain    : out    vl_logic;
        ch_gain_buf     : out    vl_logic;
        ch_gain_ldac    : out    vl_logic;
        model_sel       : out    vl_logic_vector(1 downto 0);
        ch_emit_recv_en : out    vl_logic_vector(7 downto 0);
        ch_filter_sel   : out    vl_logic;
        syn_trigger_start: out    vl_logic;
        syn_trigger_pulse: out    vl_logic;
        slot_idx        : out    vl_logic_vector(4 downto 0);
        mf_ipcm_acc_out : in     vl_logic_vector;
        mf_qpcm_acc_out : in     vl_logic_vector;
        mf_iq_read      : out    vl_logic;
        mf_choose_lb    : out    vl_logic_vector;
        mf_acc_shift    : out    vl_logic_vector;
        mf_cycle_num    : out    vl_logic_vector;
        mf_err_clr      : out    vl_logic_vector;
        mf_err          : in     vl_logic_vector;
        sync_slot       : out    vl_logic_vector(31 downto 0);
        sync_encoder1   : out    vl_logic_vector(31 downto 0);
        sync_encoder2   : out    vl_logic_vector(31 downto 0);
        iq_buf_write    : in     vl_logic_vector(15 downto 0);
        iq_buf_rst      : out    vl_logic;
        shadow_cos_sita : in     vl_logic_vector;
        shadow_sin_sita : in     vl_logic_vector;
        shadow_choose   : in     vl_logic_vector;
        shadow_read_addr: out    vl_logic_vector(15 downto 0);
        shadow_read_trigger: out    vl_logic;
        sc_status       : in     vl_logic_vector;
        sc_sin_length   : out    vl_logic_vector;
        sc_resync       : out    vl_logic;
        sc_err          : in     vl_logic;
        sc_cic_rate     : out    vl_logic_vector;
        encoder1_dir    : out    vl_logic;
        encoder1_start  : out    vl_logic;
        encoder1_div    : out    vl_logic_vector(29 downto 0);
        encoder1_cnt    : in     vl_logic_vector(31 downto 0);
        encoder2_dir    : out    vl_logic;
        encoder2_start  : out    vl_logic;
        encoder2_div    : out    vl_logic_vector(29 downto 0);
        encoder2_cnt    : in     vl_logic_vector(31 downto 0);
        reg_addr        : out    vl_logic_vector(28 downto 0);
        reg_writedata   : out    vl_logic_vector(31 downto 0);
        reg_rd_udp_mac  : out    vl_logic;
        reg_wr_udp_mac  : out    vl_logic;
        reg_rd_sc       : out    vl_logic;
        reg_wr_sc       : out    vl_logic;
        reg_rd_sdio     : out    vl_logic;
        reg_wr_sdio     : out    vl_logic;
        reg_rd_iq_buf   : out    vl_logic;
        reg_rd_shadow_sc: out    vl_logic;
        reg_wr_shadow_sc: out    vl_logic;
        reg_ready_udp_mac: in     vl_logic;
        reg_ready_sc    : in     vl_logic;
        reg_ready_sdio  : in     vl_logic;
        reg_ready_iq_buf: in     vl_logic;
        reg_ready_shadow_sc: in     vl_logic;
        reg_readdata_udp_mac: in     vl_logic_vector(31 downto 0);
        reg_readdata_sc : in     vl_logic_vector(31 downto 0);
        reg_readdata_sdio: in     vl_logic_vector(31 downto 0);
        reg_readdata_iq_buf: in     vl_logic_vector(31 downto 0);
        reg_readdata_shadow_sc: in     vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SIMULATION : constant is 1;
    attribute mti_svvh_generic_type of AW : constant is 1;
    attribute mti_svvh_generic_type of DAC_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of ADC_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of MIX_NUM : constant is 1;
    attribute mti_svvh_generic_type of FREQ_NUM : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_PACKET_TYPE : constant is 1;
    attribute mti_svvh_generic_type of sita_w : constant is 1;
end controller;
