��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�	��t�q��Tj�����E�u>�ET�Uj�a:W0�{E9�0#v��g��_e�I���7���eW�t�Z�.1`��u'�8�7p�b��I)�XO���n0����߲����7ɬpÝV�%�T�g@ ��bٺ#@���&պm/X�b��XU�PаgEn��8(�4kT���(F)C�)�@�ޑ�Um-���T�56Xj�}�ڴm�nCO�8���t7ྋ�ߧրkǎ~hc�U�.sТ���?��yk�0���)��I!��I�>��Ўru����}���T�-?�"����$$��%B��/��@� ���}y�ܞ0h㷴�<|����G�֢9���n<��|��X�?k(��x#�b&��ӽ^�,ܴ���X��jNȺx]�^r��`sNC�GVl	x<9L�_4���أ!���m�So#�r��vK|W�S�a��Ѿ�U��<����=�V ��m�r1��&�4n�>{�6���!���֎ϑ$�1pQ�I�'�<��>�N�R?E�U�e�.�\��n
���SI�q5�;���3�?�n��Fh�[*�3�`�pՔ�Ya�e~Ù?1�&�8��; �+��v���zXǡS&�p�wK��.v+E��F�-�g;^@7낄cqif��s��p,�'��L8K�^%Tp~$+4���f�����7��(�� �|6?V�I��w�n�/~�ې���׿I���z�y���h� Su�AШ�ݴ���ٔ�鑇)���K}M"oS'{iV�|�ŭ �i'T��O�͠h���c��#:�!�~>���+��RR�����g�<�A��?�P´3&��T�Oai����ND�Kv6����
f1b��m���01�ٻ&�6��'݈.B`
�q<<��Q�$i�������z���Z�K?v��?6����}�1�K�&�xj���z��-��Kn��ˤ	ڢD=z�xIc9}-�wG#��?�3�|z]��To&!��n�����6�/�{��ކ*� �m@܋��J�$����N���%g#��18ƹ����"N���~���l������Evd�!�g®���WL��H�R�`+`Tc��@�l�۵2�cSE^C8����-�U���z�3I�P=������m ����&�����e�7l��"2��Ԉ�T*��r�u�"�%����Jn;�]k�A|W�ԛ��� ���B/�+�i�	�F/���~-e�&^nfY/H���.'�|�_��0���j��"觹T~�=e�0,v<&Rĺ�@
�VV�nn�a�'�=�T_7�rT�6�	�O����v|J�x�"RBVqL�c9�a�����J��h���[�jb+�!�M^��(�R�̚�z����6�l�G�����Ztp�ǩ�L�_L��uN�%c���i	G���Ò]59��-�5/�n�ƍ�V���oWf�ؐ1K��!���o�K�C�Iv�ؿ������6�|��=�Xr��{�7?وv�_��[?��\!�+N� �x��J�$��9�*w�����Y�˗jYp��d���>}����@�������j~"R:�F5Y�}��8>�lhYD���l}챳-�J�p�	�R���\��+b�����+�URe���_����GN�sz���u�0,�P�.�ҫ�ӧ_�8�h�8{��C�1+=� �K��<���I��m�}�0V:M��*�-KS�#&��kf~a�#�]P�N�9E�'��WH�09���Yȡ���)%'$���蠼�uA.p[��wx/��@�x��-���Ó�(�9.α��#[zR�yo �m�#���S����P�|��ȍ9�T
N����_��LZ����i;��0�G���f�P7ìQr�X���L�2֎)\���q�[78���
��P�\�u��P��5�����[���^�T=� �Ֆ9�í4�0����Lrύ�f��"�0��NE����;U@A����M��٧[챬:Oh�8�$v#z/��w�z��X~��=�a�f����a�"#�ے?"f/��ߤFJ��ln�t7���
m*W^�˶�F�=�����	]�w�*R���r�RwKi���i�(HW,�=HVY"� ���P�\�X�c�Af�z^�_�-���連��b
��G�=ט��-0��(�]�V?�x�v�i�*#;���#��r���u�f�`K��AM���S���x-�}OoF�MJt�%�iu�r}@�Z#_�7�u(���"}9Ɩ�%��>'�j�$7� �N�(|�G���3�s��_QJHu���DM*?�Ygm�j�m���r0�[D�춙�,�"Є7��YI���=��,�vZܪ�A9�x%]�0n(�T=����i/�Zm�	������xt�R�W�&+<�]&�*S��;m�y-�I�_�C�-[�
��UM9ث�EH2�6ZQ���VN�$��XNPt��9��Xd�����ۿ�* ��l�E�xpG~F�A��I?�D/l�w'd�`��T�Pi�Y�@B]z7|0���)������������ �<a����x�F/ W"L�㷊!�	IA��,�7�cȥ��~��ps!;��H�qa�d��g�ox��©��锺4�i��A�Ayئ[�9�����6?�i���2F�qݫ!�@��L�B�cW��#��R����?����-��؉P�y�<^eG�C d`�#��	E��s��+��1�v����V<�8|$5�ی?��+B$�LDq��/�"v?�	�*\�����vk���&����>��M��d��~R�bl�6����2p��LǄ�5�	�>\�uzV����m�}�J"��(�R����ds ���f͵κ��6i�S/4���S����+���U6����\Ŏ�~:_O:���^��̰���P��b�5b���ſ���cn�O8dv���햓��d�[�P�������z�_�D�7p��V�x%�l����6�Y�8���'���{�_�;��5��`������Мr	O99�ߋ�=B����Kr���Vz���!�/��P��}�6*3�hcO(�Ut�צr�mv�5owpD��$���U��AT�"	�`�==�@A��|�.&�皸@�$xB��/"HI�Q|lJRccQ�&:{>�9��`�b�A��(:0U̚r���p��:�9%���7���Q�b�_h�͊I��)��Q0E~W'�������������r[��5�p�rg-T\�*6L��lfpw�̧����sJ��Ur�AE���a8A��P%���e_1���p5�����2����E)W
n��F;��7b�dGs���Cú%�`��z�#��t���֩������~%w�����=��.��(��B��������#���q�^�v�5H�ֽ�BkN�$�"^�>�؏
����*�j
�ްm�%@�~�T#�&�=�T:�9mJ�(g��B��cx5�٢�#�:��z�X�Э:�iYF�^���sޙ�i�2>wc�i�9>]kVHS"�'az ���6�y�+"��Y��T�뿥�o'}�3���lpĉ��)�l�~Fh�'���~��f���F��W��� k�u6hM��x>�N��&/0]��zn�iKCA�����l����������5F�����T︥�w�*F�ka��3�OAk��|��33ƹ��ڦi�[���P��\�;��(U�Y�=-˩?�[��t��1�_���1M���I�w�Pco�($��{$���\�^j�Tiף9:FRG�W-$��덅(���5�fy���Zf���K�,�Ba���Tɤ>��@X�	e���PL-ɒ�$I
�gM��:�㼰)�e�%"���	���T�S;J�l���T5;�ɦ@���<�e��Ʒ�=��������{���a��;acD#".g��t|�?��Z�L�}��z�K�Ǭ�����&xn������!���ޑ`@����cx�e�AhI�K�].R>.]YV-��A[��kp�·�����7n�a��2`bTf7.�d���m�1Y;���ا9O
}�Q����~�r�)Fm�)��+
���� �Pl�[(�٦0[�RA�tsģ��Srϻ�7�ՙ\16�����}5m�cể��+.=���L�#c�R���eW�`�%��vk U��pyG3g����7 �K�]��^!�Y��\�nGpVJ����U6o�2��;ƕI+(Y�`k�+G���ڤ�D+�����${S'L	��M�����Q�5�W�P�3�Vt�S�7ؠ2�����ǆ]>�l���7ΰ��P���n�'#��\8� ��vl������j
���p�!�C�-v�?�w������Rh8��u�����$�mu�Y7X�������D���gy,n��3�|����艢ސ��:c���P�M�5l�h��`r�J��ӁE�\DC#�f���OBd�!#+��t���/�Q�k �[ֻ媗xUZ��J����q������Gz��p�i���u��S�7��8���hskkp�b�ӷjpE�T��x"+��Qu2ou&�-\B�D�w��+ᠶ#9��
y�-~�@͹��~���4�_=/(2�1�S[��̡���}�cĨ���AKʔf��B�Uť;��T:�v���S�Q���O6������]<	�x����F��� �y�UM;h�$}�����B�]gSL��{�����7��.��m��~��өi:�� �P�hU��O��k�ҩR�G�T(%9T�l\\l"E�w�]��&9�;<)zkM�T�-�����k�I��s��`�cŹ)GD>��>�N�������E�K�(o���7�Oz*�3F�㹲O��F�%�ס��E��ڎ���m��==� >�>���^��M	Gt#���� ���+~"�7��wKR��t�M�����Y�-��𱇝n&����Fdh�Yt G!�<�9uSү��,�F���Nv~_��f�FT5mI5͝f���9��
M��K&'�n0ĤQAᩣ�!��xYo�B�̼ �2�2���$��'�޼�zOa-�w�c��d�o`Y�,렜x���� ��WI!\����g��mn�N�=è+' B�[gSA$$a[G��#��
ľ,�5*j,��w��2�]E��Cc5��褤"S����6�yG�uz��F�X�Q�5���f�C^�������yj��K�6�F,;K,�D�ח�½8R�l=�a�/��d
dq�D������i��R����w�{�Ji�k➂źߺ
���� ϼ�nT�[���L�)�����.��'��bDA�����d�;�u�����Hv�Zݘ�G�Q�Bv��9���D`�|8}'��j|�{}�$�P�{(*SQ��yX�~�R�?����փZ�I`ୢHL�>�
l��iS& �Xą\�0ED+��b���`X%�+�Kz��wn����%�3�D��� ~��k	��C+�`���l�m�E�8��z����S�fJ��tB�@���9���*F]!�(r�˛NQ5&�ܴ5�C�{`~��� y+�fa�@�����Se"Řko9c�9{Tv�;�v�hS���w�:����8�s	��D<E]�ְ����~��G5��邤����|�F�FL��v�P��g
�mZ���E�	gJ"O��;@�q��b=?Ł]�L�S^$ĺ(�
�3���U�
r��dc�_��tY׿[p�J$}�nnQ7��;�j��D,^�O6�k����p��$^3dց��X)F��PI�f�~P�p0F��ģ�.�T��-6.O�W�܂�Ac۟vI��ݰ�ğ�|�oƊN�%&�����w�J�H��I������&��ʯ��jm�HѬ�r��.�z��&�����P�:��*�2�����s���˨�~�N����0Ӛ��ihڳ$��fm�~HC1������̉�b�٬�f�_�Y��y�t�s���N�^(l���s���/�Ǎ�]�uV��lv��0[L*%W�5l�CQ�|��� ��Z82�C'��}��ʥr g9EK]�S�����cH�O���+��b�W�br���ƅ=��2@&���LI���W�̊	���kG�}�k����x]:;~�*d�.�PԶ;Wo��)�%Ӆ����l�Yj��Lw2��w��m��
��@�#1y����p�N9�g�)�I0����9��k5=��XsS�3�y�I1W����0	Fҍo~c�:O|�;liB�����A�.��]=�� �\�v)��Nj�ߚ|�������7U|��;9����}��`����	� �<2���I��,>\}#ʦ+�8��.d�B�mo&ڎVi�h�4e�n�j�Ϝ�i� ��(�ڦ2`t��.;Q7�Ν4�LXEO���UP��<������ö�ƞ�BUBc_7�)p�ROR�e_�g����2HF�H���deJ�J����!�=9Hq�4xt��E�	���B�5)M����WQ���Y�<��rZ�:��A�"~��Ù�SF���U�}�� L�P��@��$#�������x��Q&Ԃ�[8�p����n���>�Xt�B~C��(js����_����g6k�ז�N�(�S0�b���`����鸵��@�f����@p�FZ��P�&�J��[`��l> M&���޼�!6��i@s�x���s���=:Ub����_���WYd+L���Y��>Zq���o	sF���PZg�jD!Q���Q������[��j#������t$ż}��7C������F����6*�~V[�<���Ƶđ0̑�0{6v!���㫂�GP��Z���y����z��~!?�v{dP,����dعT�j]�V��2�ʌ�H���
@����L~zX�<&�t�CF�uF���i��&Ç���Q��L.!���c1*�>Hw�VG��,_j�2��)�QDK&HmT��ր�n�ֽɸK�{[Q���;������� X Ƕ〝��\�Jϖ��0$�+|;K[=���395K)��Oqӵp�D4�XI���*��iS�<�������r� )�tl�����D3��g�R\�4�h��ʦt�5��jPN���&��ŵ��s,�G �&84c��lDHD�`�i�o�Q"=>�`;}:�s��@�fx�@��?��d�&���כ�[��