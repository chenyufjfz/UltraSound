��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>� 0�ʪ�c�}@�+W���#��Uj��mrϐםv�����%�͂�c���&��iUd]�)Ve��,� ��$�aWg%��4�J5�W�y��(�>	_�3��_��HV�x�Y�κ͑ԧ���.��1..PeZ�9�X��W�w��K�d���Χ�f m�ԾT�P�(?���[v�|���Ma�X�Oq3��n!;���ݫyA�.� {��[P�e<Y!�5	\�ܬ�pm{#��g}�G8:M_�p=D��?������m�xs��ߒ'�yA��@'���c��Ԟ�|�=}�"�q$q�12?^G�Ԗ�⿜М��R�Q�� �¯aR�Z=�敆�d�O,t"m8n~�4nw����|6���0ʈS1��)��j�~�&��sD~�S�h�P����]�4X5+cO7�`p��p&��6>,x��4���������6,���*��-����-ֱ�1���V�����	�pi�� K]��d\I�=�5\Sv&`���T&?A[� $q�S[u�kw0�Z�j���EȪ�Q�����j҇�x� �����g���u���
����Pb��ct�$��#yE{���'\����͉�_y��̸̄�� "r)�H��O�!�3�C��=���Y�1 >뀳ITX+�Q2��短�Z�0��B��g��g0����l����.�K�R�?U�΋(O�ٹ�ӷ	�bڕ���ɰ��)w]>R4OVSn�(�L�İ�H��)e%��\N� �\���L��Qׂ&�շE8fO2	�;�����`矫��)�V�gs�T�o��fd,p�Z�/g��qW$��^VHō�`��:�<ǳ�F������N9&�s	�+��{�eh��Z� ��Z���ƴ9�Lܩ�GL_S����/h|:���ñ�*q�'J����,ާ�s�$����˜��_�-��r�	�
�0�O���x��-�Gu�</��k���	u>��L��bj���N]�E���DFF����թ����<�$E����W���c�b *0c�
��~�ｭQ�;�2�Cr؂;ѫ�����p������LʰLƆ>V�����aR�� P�QScc�sϋ�S�:�D�����������g	� �+ٷ�UG�G���1�6��ճv¿���5�4W	|���ʜm�ڋ4Ʉ�7-��XR<7
Tt�c�j6+�Pv�=o��I��� �w��z��R\*���o���MiJA�!����M��(���q0�u����7�9gġ!M����q���!�K�m�/��{��BZ���?/�P�&�yW�����k"���e�6d�'m.��8���ݲ��±a��������t�e��\l��� ��&�K�_wF�Ѭ�e��,^V���Q��/����*���3I���S�r�t\��{��ǘa���ʸo<h�Ͻ|F�0���\����ƈ���eB�L`i"g8c0�Q=�eA?�(�	띒\wԹ�{1!V��:֤����J�bT7/4��
�yz3MbkH�E*�rTk�Q<x��0��0�y�'�Y.1�8�aͻx�U>1����Y��3	���S{���`f�*=;�Jw[�01��w�X�qG���E8���(�q��Ի���0�p�pQz��҅��Q�)�AW5,[�����Н�~I��H\�	>�YS<!!���^�����+�a.���r��Oj�������y\C�ȁ���٩� �Ņ��7��35�6��jx��,�`�O:�6{����Z�n.�6K�C����- �y�7���D񭱹���|�u.��3��5���m��r�R"�o��1��_e�_UMO�{�	Zu�����.����/ՆC>oY��ZqFLnb��Yu{Z�uU?�vv);�/���A#�,��2������qD7���Y�Ѥ5y5*!��������_�AU2k�f������T������bEi���f��`<���; n�\ή����lxa�i��d}�ːKO"Lk�@�Vjja�~���b�+�s��T��`��~���I$t�kؖSq_����(�#7��5+�K]`������?�f�%����C�hvk���a,1�����ν����:���Te���+�3����>���?��Z��C��EE���+h5jjq���:r����4�k�����+��]�?m����-{�q�0v��j��Iy������pK�%���
����[y��y~ϭ	5��ِ����ٍ��}��!7h�<���F��������:���}�X�+$��̭�ۂQ�hR����K�ɩ2�]ʍ�u���r!�}P�(W�]1׳[�V��g;�L�Ԙ�H�kg����������o������3uƘ����Ŭ��)j�����%+a_������No�u>�Hg|����@����4���Й>P��e�*<�d�^�|n��`���*{��R=� 
)(�lE`��~��R�a��]G&�I�NO�;|�"*f(��xR�Dm
	|_�!�)ѭ�{�B���*Œ0m��_�y��*��H<�[�/�j�`Q��b��J�k��E��ڎs�Br|�])�~۫-;$aNؘ��z���ъ|�=y�z�v�"���߈i�c"=RŃ�$e�U�N��S�'	u�	_ D�aa+<����~U�kdjѿ�^U�"���vS^7g`��f73T�O:��kL�ȥ��wh�;e#.P�؟�p��j����
�Xf�n��%��Xik�#e+pl�������"��?���xI�`:at�!��I�wRa��������B
|�܎���>�TN��p����Z�gS�+�=�X��Rn��ς�boX�X	��/� nX�4V-j��(���?J �1��x�����/�s�,��PY�m-�C_2�^��͍�!��:�}� i)]��o����QƭY[�Ǧ��1|�צj���h���ɸ��Fgd�=xXRzz1wY�k���@6�0m�"�G�?�<7�4��bм������q��XG��M��s4��Xr�
�@:�64���ژ��Vx�<�� *K���~��Lu��-9���v�/�s<I�C@ۻ�a[�C����M*�ȹ[����8r�pκ�?>�f��a���2F�w1�/���������7{L�m�����(�XsO�'�u�5�;�H`y��^~��N_�Ӟ�|}�d�?|���@����ǋ���B�j�?��m�{TZa�d�H�o��ȍ��/X���-��(ύ2�����ي�ʃ�bM/7���&i��
P^�����P�b7��`�$G��J�煏���T��������pFShܬ�*���L����1����gƁ!^�U�d��T�l�D��