��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc��3@���;��̵*T���që �|c\
��`P��o]L̛�鿕Z[<eLl˭�W?�;���Xo����^����Z�<�F�g\CT���/4�Ǎ�@�����(�Lx)�EF}��N�QÑ�*�����Zf�ϏJV�E������V�M>؆1"��0}��{�ƽ�`G�%[�,s���>�ӹ*����ںA��j�'j��''$���F�Sy�,�v��i^ٜ��/f���.�n���WG_�kQ
-,�.UI��ۉ;��Y��ULCͷ�,lY{
��B���<�����N�CĖ�Y���3r�����M�Y���s�<��4y���k�ԁ��b������m��4愥��yF�Ls͖���2w�q�����ҶjQn�C4�Ji�t�*O+@M�Z�
��*&��S,@j�|1Nf��6�F���\Ay_AU�ǻ�yq�i����{���
m9��-&RY�l|��	˪G[k��;�*(y�M/�sI�H����J�����jf��@�J��́0�0g�vvRyZh#���������l?&e��-�8�������>
��L��9�J,�3�-bo����%�2�W+�@;�*N{���}]�z�81rJ�����!7�G����g惛��J|I11��sj�܂��҃��e��="����T�e��j��$�a�� +eǪ�
r�:��*T���r��歛}����Y�&$ ��W�E��~���]��[w~U���毀�p�ذ�S�1c�m<|]��v���"6c̄_�+I��[�3��=9�A�� t���+�7�e���\m>�f~mɳԙ�)TL'ji
x-#(��I]��ϑ g�PGrB�4�Q�.F��B�՛��L56�Y���P��R�C6��>=�u�3/u{CF ���E��s���K-w2����Ԏ�J$�
��j���2!fւ�zL$*����NR��Mc��aT-������o��(������F\D!�ࣣe,��a]Ky��n����׏������<l�]m�<H��T�X-kh2��/�$�y�K�9�7��y�.�A�A#g|�M��H��Яa/h=�׿k����X̽Ӊ�m"�6��jwl��]|Nڿ��\Ɵb�J+TIj`W+oE��1�NӖ:SZQ�Y9�ω�mC�:P�h�{�
!��'����:#v�q����~���Jz_�ȹH��ݙ�3t*���Ў��Ar&0�#v�c��Ri��%�5��%KCw6����o�P�Xѵ��FG!D1��,4<P��ɻ4d�ᥝK�;��n
��lV@�֬}�Z⡼`�!B��r�a-���Ě4Sam��R)LR>��Y�O������Y4�^0"M�Ä[�H�,��m=�(Cu"}6o�`c�`�lNe�s�T����/ٚ��T�A�~Ժ@���k�d"P+�}D�uNF���_#��,8
x��� )X�%���g���7X��#�fD���H
9�>|��
��?h�wT���z��=ti3H�ծ3��v�70����io�Yў/+��4g���`@����L��n������l`�*��������YB��ޡW�X^�u �9������5K��hNeU~��w�Y�=
�B��^�s56P��� �;)��g��6�j�i�d�%���Hr�����o�[��\��p�X�s�#��rɫvv���%�3�E����~�_�xֲЊ9}��Z�-�n@FZm�@#���@Ԥ�ɗi8�d?�p���5q�U!��Qy��s�����	�2�E+�Y�� =g�XO?I�����v�V@y|*�=Dᛏ���P��q[�P	~��Y�p���NK�1��<�yp5^V����_g}f''��?%����4O�+I:x�&��-�Z Ϻ+,��F$��j���>�:W_�8�h�li���
.�^��K��'������}6�&��#� 5yk�l�r�~M���g��4J$�M�x�v����/�ȉb.��&�"�Ī������仺��x��N	���������5��0��ϴP-�.)�9�oail3j��dݝs��_^�����3M�����Q����`n�e �9T/^9��+�$>�sJW���9�ô��v���@ǻJw^�)|-t���M��S��/�9w^�\6 ��%��8���`3�}�S��$~5�c�_5��5�J⚏	_i���\zVN7
��\���E6{!-w�^�ôtOS9�M㱴pV Ba7��<�@��5������6��[�{�珺��Lۿ�����(>� ��_0��8�dKߣ����L�|. �oˢ��P�b,U[�[�ܳ�d��Z�AB���I% /d�k���A�M��M�'��)���D@0Z��7~������Xx����|;H������Kvo�,�FO��_�D⿲��̍�&��S�yK�wn����<a/kU.icP8a`�g0�<��I�j�o�%������{(�R+V�X),�#�9~�!$�� Q/�rDűCSȣ��O�Du�h�L��E�ͬ}��MT�r`�/
�׫�E����)Q9���#��.�07=���������DG�F�
�b2�]ӧZa/�(�X�kYL$�xmw�C֣b�Y(��i�}��@����E�GF�c�/����KMӝͧ(�N�rN}��g9Hy��͉�3��y����&__��YA���Rk��02?��l�w��f�H�%�l]xW�V�ī��ld��d�S�SA��_m��J�7��g������x���;NlF#\��:��S�95%5 2}�S��n��_ӯ�h�ג���?j�D�ƉQvh���5��j�y|y�g��B@T���1[�
}����T u]��/���`ǜ�oH���w�e#�mA��s@���E����d�� Q�Jy��zG�s�J>d�� �P���1rj'Vȳ:&)�v�m�?�7�ټ��H39���s�A2�ï�R���T�>p6-