��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�7ټm�lQ�חY����C9�n9%�A�iN�k7�r���D���v�O�P�V*�d�����Ρ����Lޖb�lP|�����,yvJ�O�;Ҙ�e��< _(�����637��k�g��t�+'�����m�@��5֔�^Z�mwG3-�%Vo4x���\N�,�H�y��/
�.�S����/����Un���i �f����#��� ���IW�`���(�N�P#{_��� iOԯg!}U��(ޗ�o/��*�ӘH�|�R���϶L�VyO`ec ~����/3v`8d1���p=�b�Ir�`Q�*�����+���!�M��H�#Gk�o�{��L�7���|�f�f��с���������'��h�՛�ߊL����w`�dY�������8�c�XҮ��T�G�0�4%
^K^6#��Ǭ#���T�4����$B�>��'l�nC=�\�d$NI��Ƃ�ƪw�O647�[7ǧӗ��=�"|0��S�=7��l^l�B��n?�eI0��]
��Mb���rB�fKɆ���_[�W����˭ ��-�5�{L7�QF�U�T�cUI/ޜ$�ƤZ���{�QH+g䣙ݚ<�띯P��eFѮi�5�K�"��c!��#�����4��/Sto�nxÈ�v҆
;\�Pk�浹�g�)��1�E����ȟ ���Ө�������E�y��ͫ*�%<i�/*a$��G$��m?���kv�V�>3��Lj>���K�� �[�#�g ��de	�B���Q��ul��S[��b�KyZ>`O-Mބ..�|cN���^Ts���@�qa��l�ڰ�!�����P.[�8�.��_I9�r��Y���{��&O�0�`���=r�=S�S%���S�����S론wS c����z����u+y��_�R�Sp�v�,q7��j�;G`;(�b0���L\�6~8ӄK�SQ�Y��$�oW˳5�r��������A���צ�u�W say�ң� #]I���h��A3��Y�(��E� ���Z��P/��"�r������fQJ�?������cX踺�΅����+�F��K+�CL��i�q4S�ܡ]R"F|�ҡ,û�G��n�X������p�����	�9^_YJj�r�@ۣ)�?͈�Aߝo�E�i�ᱜy��o���C�O�;��fwe�~ЮtQ�n��3늙6�2މ��i��r�̅2��`�f0�c�&i,�(�|K#N?|�%�=��ǀ-h��֮o'F��4,�2�������9'8_1������tWD�k�5�����k��5�U�k^y�XG�4YQ�v�/��i��6ij��"H��R�|?����!Ik͖��b�"*�%���ƍ�-U���=!�zGZ�+�� eJ�8x ���}q��f�ݩ��$������S\�S&�V$?�E��S�
�D�;�"��$�R��t�!�6��:��E������T��O�-�_sP��ҝ�ZP�K�Dqj9\�� ���ъ�˭��1���-�˻J�g�\<��௼WI��%ܘ�O�����D��6;^��ߌ����I��
P��Gu�*~~~[hn���Fz�HFkf�:��{��n�=�/`�o�����)4��)���f3���.L�7���0��?�y��?�1v)���Xd����j'�2-E<6[w�&Q�����v�T��gT�s��3�C@��J��J*�H�|�z/w��t	4o�J�q��Xu��Rn����҄��GՋJ+>:�n�O�q�Ф/�^�i���>B�O�,�Fa�ѮD�^uf+2�O⍱f�e@�<ж���c�`�܉p�m4���̣��O�$9۶r㍁��̘�%��{PsX�VT�Kφ�#a����[a�f�NF׹��S,��C�dM��?�̇$��Όu�n�$���6a�A
�ɫ�@?�#��8�c�06�Q�؍�䊳m�P½�ˍ@�Ҋ22ʚ'�Yp��T1bm��/vZ�F�u�H�U�;��5=���G;�^"��o_Ћ:)fB���5��D9�L7j��f衟�_�.ޙ��k�" Y����K���}���f�d�ՈxR���wA���C0� �xX�� 1Ei_��β�Ѕ��*+ r���w5�Gy-_�t��Y�o]i�sIջw|0,�`ۚ��c���T�sJ��s���_K�x�����$",�Gla�O's�c.��Ud�CA�M&�5e��x�w�'	��;.�y�u���\f�~Ȑ��9�qO���MTb.�n��g���w8�:g��:D��A+����p�ݠc���F�a�Ԍ�G�IT�h�([�X�PD4�	W?������͠��jEq��KZ�B�?,'����	��c;��e*��* M��8R+4|�����O7��9�hki����4��}��,Y�D�N�c�������O��;���Gc/XvH��	�d��K�'�aϡ�X��tFTS�䰎4Rv�7��RN|�{W	[eƹ˗I���
�J������P&��-�\��	r�L'��uil���6����ݩ�_j���C #j������h��1^Gw<���<�%z�9ĳ��o���kմa4�"���c��oﴲ�����d�G���q��ߊ"H����{1��f���7\��{!���h����,E�	�5v`D5m�CM*O �����uRM&�8�olX�6Q�p����q�y�+�7�pE�C@�w�?c=��� D_�բi��wL�)��x��,a��G*�m���T�	�_�D���B(��,�J�|�k0\i���7|�[��jjP�è�}�<*�Y���~ �b���:���{VL�.�����8��uu��v�����9�qcg�k�