��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P	����6��<����`V:�Ufv#�խ����!��O���$�opB����n����\5��<`dQ!1O�VK3.u��q�Fy��g|l�RQ̒�jv�
3�-U����X�A���G@�B΄6������{$:@�>��*(E��¶�����u(�,&�P9��3D��2T�v������S����Z�������hku�á����>�����d�rI��e�	�5�I7#�v�E\$��Pť��7�su
����GQ�%����c�Қp.P��r,����k�-֧���K4�q�0��������A�����Ղ"/y"���]�j����U��6����scS��$Q�{h5}q.1�����:��B3��ʦ�e0%�5�Voݫ�w'�!'�;<�u~&���L�U7�u���H�;΄�|*iN�T�j
&��ވ����z[C�J�V\Nu	�����1�+�TfN�M�7ϑ-P�y�R��z�L4}2����B�L��$����d�R��O�зs�'
2�N�K���Y��3gg�{�ԗ�����S��R��i���~ؙ?)��or��$ĝO�7������0��u�������j��.)_�N�ޘ�Ir'=`׋G�+6�1��柕�FO�hQk�Vp�T�s�=[���=��_y�ʒ>$��fcn�n�:l�Q�+ũ5]4l��Y������룱}·�0AOV�x��0�+a�n��z��Q��X�7㰺ߋ�G���Yc��*��~�!2�����RJ$��F<#L��tS���#��k]���
ѱTm�����k*��3ӳ��qqd��)��k���U4�Q�Ҿ��'԰��c�"���$��>tV�m����� ����`u�PX��n�F] ���3�]��������F��ޑ[xp���$�����.�0�wbw��0��Ц1���
��K�oN"X���`�4 T����]@����38��jwN ��9�jW3� ���t��5���1>۟�������ʓT�o[�tƦ��)�4�.����a*̆����
�앗���K+�I��P�e��SR��g�� )pn� Q�_�֚f�����X��q^;�=�4�Y�e���w��K>�#iD�_Ø�
z���ӧ�;̋����> ��+�R6z�M�����q�(���3��&�U,��?�P[��!�m�0h.3��ݙ���Gd�(�S`.�K�.�k@�,�ܝ��5�y�v�/	UH5�E�H��	8���\;$�Έ^��<P7&i�w�ދ�|�P�
��]ڟ-��]f�q\ey��&9@=U��K�y�#�Gh����S�5��`!F�J���yM�K��{�>�S���<`�{�|n��_iˍ���7-�G����� �?�$�P��A?,s=b��L��I�"G�'u}���o������X�}�iS���E�$�d2DY}�j_H�1��O�0i���GN�H6���!5��8;GG?�D�p�:�]@�8�,a��p ��ztB�� �����&��op��*6�gd`dV,���`'���CT,�!Oѵ<puF�~<ѹ���5Ԭ1"���{á��'�C�Q���kބ�c@C�^�m�S�ؒUM����~��ٳƭ�V�3��?����G����IC ��F�=���0�=��̓*�E��4�檧4l��������R͜Y:z����H; z�r�KP%�P�t1x�}�~pA�,;I�F(�V�J�6�{�!.��9���d�Pp��L'Z��V���R�����*	�ؘ��%�Y�Gֳ>:�E�X�*J���lѮ�9���4�g>��z�Gk�н���E��c򭹽�b�_��^�a�#lǙF�S
�.<&�)[���΢��f��)���ś�ς ��>��*���=�0��ZD�ґ?�.�4���J�B�)���;+Ev��ݖ%B��K�Pϡ��	����I��^#�!"b�T��E74J���"�WCE:ۯf�A0�)X�|�&�ں�� L��2��"�T����:��0�b}@������w@
�9��"%R�!��q;��g6�h���~���=�u���.�y��	w!">��O�fLc١'0�O���軴�3�E��H�T`��l,���kLt�'�+Z���f���t�w��7�v��i���TW��/�ezL�s��Qk�(�f��4a����ӱ��ޒM�����qq��+݃ϭ�H��!���o�}���H�׉�]mx�E������1{E�GҤ0R���1�OϝCM׉f���4�Y���~�����Kƀ���Q�����`W!".��H�0c��;�ŉSNs���a�J��?��O��g�w���LGe�a�g����]�JPA���u���cOf�ؒ�����GT�y�bL�Hj�ְ����;ug�m�`��L{S5ט�� ǃ���u<mHZ�L�H�l�H��=�}�&ZQ�y��oTA���W`��VU��;�n=ݐ��>�g	��;T�D�f�\�G#�r�FH>+��*�Kmz<f�; ���[�%e��K��5��q���E�>��=�E�&��U�<�=q�Ab7Xǟq��l_��� ��� 3֭5�r�:����|dn�Μ�M"���&91�Ԗ|�b+8n�.{n�jR�B�#����e�b�������7_�M��{�~���_�'@�Ca ֛�A�Kw"8�6��':>s��А�N6M_��x�e�t#=n��F�L9/�J���E+��w���*�-ȗ���.��r���]�U��-F;x��F�s��MR_Yz�er�����xe��_�&���Oi���I���T��v�S4*�~��2[ko2��+^�!�]d6���\*N��'�Njf�o�S�*b���W��x�P��~��Ĥ��/��SL�bX�)���BU��C�Ĳ39ej�}��`х��˧L.#�ٻ2_���{�7��E���:zЩ�
r�b����!�����Uo�<Gñf�135�5w��1�:Х2���������#;��kD���>	ƥfC}2D�M�ѻ/��Z��.=�ٕ�S,n�f�7����qq\���:z��'B[��T�5����nЈށ��wγ�K��H��M�7�pw|�D0m3��Ȭ�����C���G̤�=b��E<'#�����݃X^,�G��������ۖ0f�QJ�&Y�'�~�Ti���w����H -�%gÎ��n��c_���e��ٍz	J03��꿑MD/Z�M��6�v�����ܖ��MóMP���q��*
1�׷g���)v�6
*�C��M����F$[�R{P�n�_����7��q��DI����י����G#gU��?NtI����<b�Z'wDV{(�R0�o4̯<m숢Imb�(	[}Y��%�*���e��'�d���^�g��b3�C56A�C��ŧ�����ӣ�p@V�^���[h�����jK11D�L�^4�����G�y�51��B�y$�"�#����{��G��[������J*/"\���Qڈ�G!:m���)d�|Ĕ�I�*��o4��b�����CM3��~��m��5(��[�a}?^�aӭ�ǹv,GQ�*4	�ōf��\uU*����u�?4�e�e��$
��v�Z,����3���Q��˧H%_9�K��
�3{AĲR�^,=)�e��v,��ji{1'�9�wfw�������W�檼9�|
g���g�y�V�5�M�`�̭��`�z/g�`6�I����8��j���)���ڵ�B���.�����1����x�i�׀���42�ڬ~�t�W���;@������5i�K�a5U^0���N���y���G��r���\Շ��#ī~o�DM�t��;��N�pK�s�rf�ES=��n�#^�u��J�>Ƞ��؆�E�����+�j�ݷC����ʄ��-���w������0���d����1=�Z���E
�0j�(lS��%{#�q�[`w��H����n���	����ctGy�Z܄�>j�:/|ބP���� ?í���Q?T�C/flGx���t�NZ�|Γ��[�]sHv�.��_�2�J���
a�څ��F������{"�5� ��M�5��Bl��7��PRe��j?^;�*~��-J�K�J6O�f��c3U��Y[��d��i�u҃$>S�ΐ�eS��A���7�g��v�!8(sC��|Ն(��a���ꃌ]s<��#ؓ2��Ex�|MB�0���f�
�kP�i�,�_�0g?��%����ɓ����?�9����M`v�J8����j��r��K���2_�ېxǘS:d���m$|���}�}���ũ��YbǲV]��X`�_w(~���L���\�9��N�ܬ�P9\���Ε�����oYL_rv�8�H��*�x$�|B�\K�a9�&:�p�$!�,S����Z��_�מ Z��1��۹n���.!���msM�a��F�"?�L���5Y2˅����j}M�Ի��]��4�1��K#N<:���ji�&�ת��IM�k��d�>�-v�d냡�����˱�0���N�����<�|aJn-��jE�g�"��A	��>�HXs/���h"����c�9�R������ڟ�r�*��j��> e�Q+g�-�+�d�Ģ�",�j����K�G�-��,!I�f �j�_X�n�v�����J�PXX��u2��
�j�~�e���T�~�C�M�A����1p�W��.��t�C���o�[���OB~:��;oD�,F�l c��k�j��*,9���
��R(�W�^Ң��Sb�(�Q�UF(o�Z���=�j�2@H���N&'hl�}�F�O��e��$��hQB�Z��r������Ȑ�v�+J��������ؕ�+���oR�ڡ�>�f�pÈ���y({->@ۓR��r����2�{cz9��i���,-5���:Ěc��D��M�H]i���?7��mHh��W�C,zd��ϐ���3�|��5���
l=�p�q+xv/��RZ5�wk�Η.��a�A�/���Ѭ����t�*����>`����4�єw�灤�ь�CSe>�&{���:f�:� �햚ʱ�7,�m��}�8��c�B��]�g��{p���Ӗ:�ܾ��ل{ߖ �K_vg��Eu.��N�.�g ܪFtý���a�z'Y��I;��е�ە����#�@��㫢��`��\�ZzlQ ����i
`f �ˈ���k� 8Z����!o����x_��GJ�����jW����I��R�k�a�-׮� ��������	�"p�&�~�EF�%S�8W�����-qJ�kKk	���w"W+�i�0��ا��R�0i�V&�f��-��}����#���4�\��?"f!N�\�����R�[����*fF�����j�.�m�t�G
����?ۥ�O��z��茁�����T�>� Ά*���09�wF�4�Op��>z�h���Ě��d�����w�ػ̔v��Y?�93�7�Œ��K����LR@a�u'o�����uLI�Ć\�����l���Q��H $_��Ѡ�\9��%���}����V��H�F�c����x����wiwQ�z�p%AZ���g��4�����B.��{Y.�J�4���3���B��#脪l��k6�\�<�(���X<(�>��'K��':/)[{�&����_�qa�����5��M�<r`�Ή���g��mO��^�q:���A^|R�����
{,EI��+�\q�/b>p�ม�xE�8�9kQJd-[׻�lHg���Ct�B ��Ɣ�B×kî���_x�a<?	�K:}�Z����.�������Ű�O��r�����g5ҁ�!E.��j�~405�M����2Э���r�T�[;�����xb�l!h om�wCbۗs��$��������Ca�JӡU)s,�Xh���~Kv����dk�O�0�O8��[�jO?|��9�l�2�02�~t%��1�� u��5��~e㸐�׾��߲��#���n[L!������B��	;lU���>`�q�b��,�� �vm{��R�ZL�$@��e��@1��h�b��`G�0�=��+�F�]�@��Dq'�bՉT ����`�t�W>
_3fSo$��y��! 'jh�D�{��?��?�+�et����p�@e�*3�{�J|ih��$�\���[\��C�)-.y���@v���vW�Z��Ȑ�m�)u�Ǻ�Z���l��ng(��zS�W�ϐ�W�U�i�,4p�qGv�B��#�<��u�a~�����@JX�T�렮�rE"��`XO��C���n$n