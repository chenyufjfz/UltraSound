��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��l_����b�-Vx�X�w���<��l�~�s,�ǟ.HIpd"q��o=�JQpk�e�A�:�G�bV�Q�O �R������U~g<3���%����Z.���a��L��$�E>#�V��1u�Aѽ��)�G��*��jfMـNk�=�<�✈%	?$���-��束�I�3Frf��k�|u�����0΋ʗÛetB��>"�Qq·��ar��ھDB���֪��@��)盖��=���T�w$����W�Z�B��A����I�Z��M�&�
��94ݟ-7Sg��I�~����s�k	*x�P}6��+����d`u�x�	e�R� E�����Z��'�^,��P�]�7%n��(�N����Fl� w�ۜ���0����I
Us��)�C�Ld-���94�`D���Q��4%b�����v�p����e��������\�������q3��2J��	�x&��%*��h�ofOy	E4���-z��I�}dDI�Q�O�,7�.V�P�	��}�.���}�f� ��P�}ri��x'x@ɐ��洳���;8>p�}6��,���_644����K�o�':c<��ù�!c�|����H(��K$�$樯���A���Y�W��2ߩ�d������P8rW�A��s;�wߩ�N�o��?Dp���w��PY�A�-���S=�|��=���q�^d�VU	(B�5�2��u��%�a���hs��_ߗ��n��45�ڶ�n�8�)Q_�e������/m�ܺ��K��(������| ��et�iF=���f��o}�8D�+i��G�:��P�,��^êձ�;�@9]m^��ߧ).�>����k�
wȮU�Z)j\(4���K���H	�	53���sw ���Z�&,�PU���vy�ض2N �dk�G�@���JDO�c�u�)�<�?��x΍x�ƍg���|��[�4�w~��}OƗ��ƕ���ReV�D�ZS0Y�m��gt�0�wġ
v���C��۠;puJ/>6���_�zܝ��uPŠhb���Fh��LSc�<yz�0��Բ��)�X���k�^O��m�"��0�5i&���X�[���Z���z�D4�;���u����(|t��u@9�8=JH@e �Q�-\���<�.���"���=�Z�A���|�bC�4٭C �֔%"�{�ɉ�4:S1� ��Wr_����0����$|I�KF��h��>��26.Y�e��8۷��|̈n�P)3�x�f����_�ෙ�	�Ql� lbt���%r+Cz�k2ɽ�bT� �hd���nM�.�+h�A��������������C�죭���?��O��:]����뻏}�k'0�L_*�~l�s]�{3�.z����[���9[���p�}��
��f�^t�r�i�B�FYro�����h��Gs���O�;Y�GK>I�
�Хp4��(���{c�ߍ�T%�b�̀�"���&NG��= .���(e��I���M�Ɯ���R�E~-�ʙ��zq�[WQ��#�2F(<��
�C���!ω��j�xZLE"1�U�{�A)�6c|��QyE:�䏓q�	Ʌsd1����7Lz�������<�6o�{͛{����D,=X˱Ą��VC�*=��[W��ݗ�Һ#����~���.cx�Clu�$!�k2�4�3�mI�^�����������f���o�_!��j����bz�3���
t�ڒ.y����x ���.�b�����2Ty���m<V�q�{�;Fp�i3���Lb�����R48�"M�|0�}rnA"&{Y�"�a�t��wjD(��b}>ς͂�JEf�z��f�|�����SyM�Uo�:8�3m� ����u��I�uf	7Z��1�xӹ�\�/kt_vj�DZ��G�=_�r�D��[��ye0dl|F�\ʾ�$r�Cv4���CC�%�똓|��2V�\<:���\���$�h�2)Z�2ݿ|r���G�^-e��|�
9J��3����(���>��%��4n(⬸S��	�{X�k�����T8����k7�I�$���w-K��M��N��t�gCzt"��axő���c�{��f
�$��0^E6���c��ǡ��ߑS��m��p=���S3X��=!�!�7L��R6F�!8h��*��nm�A9�&�ǿ����1�
�B(�"�e�)'
�Ũ����,���tWu�n0o:F�s���[��ɾ���X�}	8/L���@�����N�
��\�)���,J*��=笶�2��������	�J��Ĳ�����N'�w��Lh<�1e�/����𳎞}1��H�'T�_c�V�$�����YH�&{]�4�q)|L��ߐF��Id׍�@�~V�1\K����p�2��7�W�}�-
�ⶩ�}u��AFa5�N�FQ���#H�4���#*�Gf#]�
�*Yշ4J����I}J� ��K1�a��+K��>v�6�V�F)��nb�+���q�@��fn��VŇ��?�E�/$U�zuȜ@_�����Ԛ!��s� �j�?砒c�<�nj�E��9+U8�$��s��m�������uTp6MU
#�!��tqśε��O^��\�I@�r�O�|�$�1��d����R��W�Ji��Ň�љ57�q,�:�t7[T�K��1R�tٟ�A�r9�ZQ�=Dk����i��:ۇ��K:J���G�-���`N�ي�<b�����~(�!Y@����m.-q���=�qL���|R�{=#�h�9�A���N��SpQ�4�;�.�q�����n���&��V�C��5����뻃�Tbvt���?�8-��3¬��J=��{���dE�HA��|
g���q�-�h��.��al����j}buL\yD%R��0��ѡ���kdZ�3L��D K�� ?O�=N�*
]&B1"ˇŉ��sPJ��"LK�*���04��&�]�R�/����Z�H� ͻ{CT�Һ��*x����?�	�:ȶ��2с����4��@�`��0��ޖ�X�1Ui�y�^]�>�yG��'�z�B���;߱��{`��2�ׁh�J|�jrn�H�{1�F�}FϏ�_ErxBP~��Dr�� Z�V��t,<���9A���\������k3s��h��K5��B�������w�:sT3<�I�?�4�sdP:.���K�fJ���*S�g}"���g߇��P*"�%s�ctW����WjZ9a�Kz�:�w�1����u����s���T�>�l�V�z͸���Nʱ}x�`���I��J5��%��7�E�ހ��?�0�����Rn�0���Y&+�7�>px��	�-}�$�N9���jT'\���P֤����3���C�|퀢X`k���j+k
�D��r�i#�w��i�wy�б�dŎHd� ��骟�b[oҡ3/�p�^Z����t��޾���~��"!�� <D<L\mu��@P¨�B���M���~��q�����
мT�����9�rY���n�+�{L焯K6�z�N�R)^
�"��h�g#p}�[��K؞<O�/^�
�Ԅ0��Q�d�a�9�����rrb��tH�yP_�+�5�@��y��� ��V"��d5�����Ư�6���Q`���6�g4�~����J����4�W!��̵a��Gb�I
��WW�s��D*�I�`�j��[�~�����`�|}�jG?�b�G����0��7I7�R��6�5���ޛf{�.��l2�=���f�%�/������7�@g�u�T��{�����@k�N�IϾ��I#�a|}W���(s�嵆l��C�\�'Y��cQ@
U]'���m3(<U�!:���kH[�K���"��o�{j+X�C���&��Ds��ĩ�!�I���	í\��s���aJC%X�[t1!�p���y�� M]L��
��j�o�hb���O����lP�WX��jAc��-r3�aJ�@mda��]���u1ꈭ���*a����[��4���8�r}�j�V@3]���%�"&����6�+�t�O����e/tz���jj�0��a�k�x�rS��Ek��rA�e�7�_��f~!y��#��{��k�KR_����(�	���8<^�A���a=u`���1e:}�Ҩ@�+BW8��p�1�J��Q��<$^Ar
�� i4�WS�h4����t��\Qpp���\uP��#旴L�Nq˲)7�r.�f�ks��KXJ���'B��p�0�\E^�-��԰k���)WW	5۫Z���8�cjn8!58P�Ø�{G����I_�T���2���i����#EZ� �ޜ����|� ����FpZ=o��H�Թ���y��c��{�R��}u��,I�\v���L~L����8v��ߌ�H��P��B���q�/�$��