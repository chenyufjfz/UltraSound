library verilog;
use verilog.vl_types.all;
entity ether2 is
    port(
        address         : in     vl_logic_vector(7 downto 0);
        clk             : in     vl_logic;
        ena_10          : out    vl_logic;
        eth_mode        : out    vl_logic;
        ff_rx_a_empty   : out    vl_logic;
        ff_rx_a_full    : out    vl_logic;
        ff_rx_clk       : in     vl_logic;
        ff_rx_data      : out    vl_logic_vector(7 downto 0);
        ff_rx_dsav      : out    vl_logic;
        ff_rx_dval      : out    vl_logic;
        ff_rx_eop       : out    vl_logic;
        ff_rx_rdy       : in     vl_logic;
        ff_rx_sop       : out    vl_logic;
        ff_tx_a_empty   : out    vl_logic;
        ff_tx_a_full    : out    vl_logic;
        ff_tx_clk       : in     vl_logic;
        ff_tx_crc_fwd   : in     vl_logic;
        ff_tx_data      : in     vl_logic_vector(7 downto 0);
        ff_tx_eop       : in     vl_logic;
        ff_tx_err       : in     vl_logic;
        ff_tx_rdy       : out    vl_logic;
        ff_tx_septy     : out    vl_logic;
        ff_tx_sop       : in     vl_logic;
        ff_tx_wren      : in     vl_logic;
        read            : in     vl_logic;
        readdata        : out    vl_logic_vector(31 downto 0);
        reset           : in     vl_logic;
        rgmii_in        : in     vl_logic_vector(3 downto 0);
        rgmii_out       : out    vl_logic_vector(3 downto 0);
        rx_clk          : in     vl_logic;
        rx_control      : in     vl_logic;
        rx_err          : out    vl_logic_vector(5 downto 0);
        rx_err_stat     : out    vl_logic_vector(17 downto 0);
        rx_frm_type     : out    vl_logic_vector(3 downto 0);
        set_10          : in     vl_logic;
        set_1000        : in     vl_logic;
        tx_clk          : in     vl_logic;
        tx_control      : out    vl_logic;
        tx_ff_uflow     : out    vl_logic;
        waitrequest     : out    vl_logic;
        write           : in     vl_logic;
        writedata       : in     vl_logic_vector(31 downto 0)
    );
end ether2;
