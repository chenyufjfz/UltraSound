// megafunction wizard: %RAM: 2-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram 

// ============================================================
// File Name: gpram.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.1 Build 243 01/31/2013 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module rowo_dpram (
	data,
	rdaddress,
	rden,
	rdclock,
	wraddress,
	wrclock,
	wren,
	q);

parameter rdw = 32; // number of bits in read address-bus
parameter raw = 8;  // number of bits in read data-bus
parameter wdw = 32; // number of bits in read data-bus
parameter wsize = 1<<raw;        // number of words in memory
parameter pipeline=1;           //output register, pipeline=2
//parameter SIMULATION = 1;
localparam waw = (wdw > rdw) ? raw - $clog2(wdw/rdw) : raw + $clog2(rdw/wdw);

	input	[wdw-1:0]  data;
	input	[raw-1:0]  rdaddress;
	input   rden;
	input	  rdclock;
	input	[waw-1:0]  wraddress;
	input	  wrclock;
	input	  wren;
	output	[rdw-1:0]  q;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  wrclock;
	tri0	  wren;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [rdw-1:0] sub_wire0;
	wire [rdw-1:0] q = sub_wire0[rdw-1:0];

generate
/*
if (SIMULATION) begin : SIM_RAM
    reg [rdw-1:0] mem [wsize -1:0]; // instantiate memory
	reg [raw-1:0] ra;                 // register read address

	// read operation
	always @(posedge rdclock)
	    ra <= #1 rdaddress;
	    
	// write operation
	always @(posedge wrclock)
	if (wren)
		mem[wraddress] <= #1 data;
		    
    reg [dw-1:0] sub_wire1;
    always @(posedge rdclock)
	    sub_wire1 <= #1 mem[ra];

assign sub_wire0 = (pipeline==2) ? sub_wire1 : mem[ra];
end
else*/
if (pipeline==2)
begin
	altsyncram	altsyncram_component (
				.address_a (wraddress),
				.clock0 (wrclock),
				.data_a (data),
				.wren_a (wren),
				.address_b (rdaddress),
				.clock1 (rdclock),
				.q_b (sub_wire0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.addressstall_a (1'b0),
				.addressstall_b (!rden),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b ({rdw{1'b1}}),
				.eccstatus (),
				.q_a (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));
	defparam
		altsyncram_component.address_aclr_b = "NONE",
		altsyncram_component.address_reg_b = "CLOCK1",
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_input_b = "BYPASS",
		altsyncram_component.clock_enable_output_b = "BYPASS",
		altsyncram_component.intended_device_family = "Cyclone IV E",
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = 1 << waw,
		altsyncram_component.numwords_b = 1 << raw,
		altsyncram_component.operation_mode = "DUAL_PORT",
		altsyncram_component.outdata_aclr_b = "NONE",
		altsyncram_component.outdata_reg_b = "CLOCK1",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.widthad_a = waw,
		altsyncram_component.widthad_b = raw,
		altsyncram_component.width_a = wdw,
		altsyncram_component.width_b = rdw,
		altsyncram_component.width_byteena_a = 1;
end
else begin
	altsyncram	altsyncram_component (
				.address_a (wraddress),
				.clock0 (wrclock),
				.data_a (data),
				.wren_a (wren),
				.address_b (rdaddress),
				.clock1 (rdclock),
				.q_b (sub_wire0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.addressstall_a (1'b0),
				.addressstall_b (!rden),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b ({rdw{1'b1}}),
				.eccstatus (),
				.q_a (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));
	defparam
		altsyncram_component.address_aclr_b = "NONE",
		altsyncram_component.address_reg_b = "CLOCK1",
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_input_b = "BYPASS",
		altsyncram_component.clock_enable_output_b = "BYPASS",
		altsyncram_component.intended_device_family = "Cyclone IV E",
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = 1 << waw,
		altsyncram_component.numwords_b = 1 << raw,
		altsyncram_component.operation_mode = "DUAL_PORT",
		altsyncram_component.outdata_aclr_b = "NONE",
		altsyncram_component.outdata_reg_b = "UNREGISTERED",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.widthad_a = waw,
		altsyncram_component.widthad_b = raw,
		altsyncram_component.width_a = wdw,
		altsyncram_component.width_b = rdw,
		altsyncram_component.width_byteena_a = 1;
end
endgenerate
endmodule
